THERMO ALL
   300.000  1000.000  5000.000
H                 L 6/94H   1    0    0    0G   200.000  6000.00  1000.00      1
 0.25000000E+01 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
 0.25473660E+05-0.44668285E+00 0.25000000E+01 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00 0.25473660E+05-0.44668285E+00 0.26219035E+05    4
H2                TPIS78H   2    0    0    0G   200.000  6000.00  1000.00      1
 2.93286575E+00 8.26608026E-04-1.46402364E-07 1.54100414E-11-6.88804800E-16    2
-8.13065581E+02-1.02432865E+00 2.34433112E+00 7.98052075E-03-1.94781510E-05    3
 2.01572094E-08-7.37611761E-12-9.17935173E+02 6.83010238E-01 0.00000000E+00    4
O                 L 1/90O   1    0    0    0G   200.000  6000.00  1000.00      1
 2.54363697E+00-2.73162486E-05-4.19029520E-09 4.95481845E-12-4.79553694E-16    2
 2.92260120E+04 4.92229457E+00 3.16826710E+00-3.27931884E-03 6.64306396E-06    3
-6.12806624E-09 2.11265971E-12 2.91222592E+04 2.05193346E+00 2.99687009E+04    4
O2                RUS 89O   2    0    0    0G   200.000  6000.00  1000.00      1
 3.66096065E+00 6.56365811E-04-1.41149627E-07 2.05797935E-11-1.29913436E-15    2
-1.21597718E+03 3.41536279E+00 3.78245636E+00-2.99673416E-03 9.84730201E-06    3
-9.68129509E-09 3.24372837E-12-1.06394356E+03 3.65767573E+00 0.00000000E+00    4
OH                IU3/03O   1 H  1    0    0G   200.000  6000.00  1000.00      1
 2.83853033E+00 1.10741289E-03-2.94000209E-07 4.20698729E-11-2.42289890E-15    2
 3.69780808E+03 5.84494652E+00 3.99198424E+00-2.40106655E-03 4.61664033E-06    3
-3.87916306E-09 1.36319502E-12 3.36889836E+03-1.03998477E-01 4.48613328E+03    4
OH*               121286O   1H   1          G  0300.00   5000.00  1000.00      1
 0.02882730E+02 0.10139743E-02-0.02276877E-05 0.02174683E-09-0.05126305E-14    2
 5.02650000E+04 0.05595712E+02 0.03637266E+02 0.01850910E-02-0.16761646E-05    3
 0.02387202E-07-0.08431442E-11 5.00213000E+04 0.13588605E+01                   4
H2O               L 5/89H   2 O  1    0    0G   200.000  6000.00  1000.00      1
 0.26770389E+01 0.29731816E-02-0.77376889E-06 0.94433514E-10-0.42689991E-14    2
-0.29885894E+05 0.68825500E+01 0.41986352E+01-0.20364017E-02 0.65203416E-05    3
-0.54879269E-08 0.17719680E-11-0.30293726E+05-0.84900901E+00-0.29084817E+05    4
N2                G 8/02N   2    0    0    0G   200.000  6000.00  1000.00      1
 2.95257637E+00 1.39690040E-03-4.92631603E-07 7.86010195E-11-4.60755204E-15    2
-9.23948688E+02 5.87188762E+00 3.53100528E+00-1.23660988E-04-5.02999433E-07    3
 2.43530612E-09-1.40881235E-12-1.04697628E+03 2.96747038E+00 0.00000000E+00    4
HO2               T 1/09H   1O   2    0    0G   200.000  5000.00  1000.00      1
 4.17228741E+00 1.88117627E-03-3.46277286E-07 1.94657549E-11 1.76256905E-16    2
 3.10206839E+01 2.95767672E+00 4.30179807E+00-4.74912097E-03 2.11582905E-05    3
-2.42763914E-08 9.29225225E-12 2.64018485E+02 3.71666220E+00 1.47886045E+03    4
H2O2              T 8/03H   2O   2    0    0G   200.000  6000.00  1000.00      1
 4.57977305E+00 4.05326003E-03-1.29844730E-06 1.98211400E-10-1.13968792E-14    2
-1.80071775E+04 6.64970694E-01 4.31515149E+00-8.47390622E-04 1.76404323E-05    3
-2.26762944E-08 9.08950158E-12-1.77067437E+04 3.27373319E+00-1.63425145E+04    4
AR                G 5/97AR  1  0    0      0G   200.000  6000.00  1000.00      1
 2.50000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-7.45375000E+02 4.37967491E+00 2.50000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-7.45375000E+02 4.37967491E+00 0.00000000E+00    4
CH2O              T 5/11H   2C   1O   1    0G   200.000  6000.00  1000.00      1
 3.16952665E+00 6.19320560E-03-2.25056366E-06 3.65975660E-10-2.20149458E-14    2
-1.45486831E+04 6.04207898E+00 4.79372312E+00-9.90833322E-03 3.73219990E-05    3
-3.79285237E-08 1.31772641E-11-1.43791953E+04 6.02798058E-01-1.31293365E+04    4
CO                RUS 79C   1O   1    0    0G   200.000  6000.00  1000.00      1
 0.30484859E+01 0.13517281E-02-0.48579405E-06 0.78853644E-10-0.46980746E-14    2
-0.14266117E+05 0.60170977E+01 0.35795335E+01-0.61035369E-03 0.10168143E-05    3
 0.90700586E-09-0.90442449E-12-0.14344086E+05 0.35084093E+01-0.13293628E+05    4
CO2               L 7/88C   1O   2    0    0G   200.000  6000.00  1000.00      1
 0.46365111E+01 0.27414569E-02-0.99589759E-06 0.16038666E-09-0.91619857E-14    2
-0.49024904E+05-0.19348955E+01 0.23568130E+01 0.89841299E-02-0.71220632E-05    3
 0.24573008E-08-0.14288548E-12-0.48371971E+05 0.99009035E+01-0.47328105E+05    4
HCO               T 5/03C  1 H  1 O  1    0 G   200.000  6000.00  1000.00      1
 3.92001542E+00 2.52279324E-03-6.71004164E-07 1.05615948E-10-7.43798261E-15    2
 3.65342928E+03 3.58077056E+00 4.23754610E+00-3.32075257E-03 1.40030264E-05    3
-1.34239995E-08 4.37416208E-12 3.87241185E+03 3.30834869E+00 5.08749163E+03    4
HO2CHO     6/26/95 THERMC   1H   2O   3    0G   300.000  5000.000 1378.00      1
 9.87503878E+00 4.64663708E-03-1.67230522E-06 2.68624413E-10-1.59595232E-14    2
-3.80502496E+04-2.24939155E+01 2.42464726E+00 2.19706380E-02-1.68705546E-05    3
 6.25612194E-09-9.11645843E-13-3.54828006E+04 1.75027796E+01                   4
O2CHO      6/26/95 THERMC   1H   1O   3    0G   300.000  5000.000 1368.00      1
 7.24075139E+00 4.63312951E-03-1.63693995E-06 2.59706693E-10-1.52964699E-14    2
-1.87027618E+04-6.49547212E+00 3.96059309E+00 1.06002279E-02-5.25713351E-06    3
 1.01716726E-09-2.87487602E-14-1.73599383E+04 1.17807483E+01                   4
HOCHO             L 8/88H   2C   1O   2    0G   200.000  6000.00  1000.00      1
 0.46138316E+01 0.64496364E-02-0.22908251E-05 0.36716047E-09-0.21873675E-13    2
-0.47514850E+05 0.84788383E+00 0.38983616E+01-0.35587795E-02 0.35520538E-04    3
-0.43849959E-07 0.17107769E-10-0.46770609E+05 0.73495397E+01-0.45531246E+05    4
HOCO              T05/06H  1 C  1 O  2    0 G   200.000  6000.00   1000.00     1
 5.39206152E+00 4.11221455E-03-1.48194900E-06 2.39875460E-10-1.43903104E-14    2
-2.38606717E+04-2.23529091E+00 2.92207919E+00 7.62453859E-03 3.29884437E-06    3
-1.07135205E-08 5.11587057E-12-2.30281524E+04 1.12925886E+01-2.18076591E+04    4
OCHO              ATCT/AC  1 O  2 H  1    0 G   200.000  6000.000 1000.00      1
 4.14394211E+00 5.59738818E-03-1.99794019E-06 3.16179193E-10-1.85614483E-14    2
-1.72459887E+04 5.07778617E+00 4.68825921E+00-4.14871834E-03 2.55066010E-05    3
-2.84473900E-08 1.04422559E-11-1.69867041E+04 4.28426480E+00-1.55992356E+04    4
HOCH2O2H   4/ 9/98 THERMC   1H   4O   3    0G   300.000  5000.000 1422.000     1
 1.16303827E+01 7.15133688E-03-2.39035030E-06 3.65772791E-10-2.10199524E-14    2
-4.31079242E+04-3.24276725E+01 1.85716693E+00 3.23153132E-02-2.69928902E-05    3
 1.11694484E-08-1.81284103E-12-4.00314471E+04 1.90917729E+01                   4
HOCH2O2    4/ 9/98 THERMC   1H   3O   3    0G   300.000  5000.000 1412.000     1
 9.04545938E+00 7.15223373E-03-2.37005676E-06 3.60083481E-10-2.05750228E-14    2
-2.49414886E+04-1.74210530E+01 2.85441621E+00 2.33663535E-02-1.88115990E-05    3
 7.96709515E-09-1.36346618E-12-2.29866196E+04 1.51730565E+01                   4
OCH2O2H    4/ 9/98 THERMC   1H   3O   3    0G   300.000  5000.000 1420.000     1
 1.15398246E+01 5.34291432E-03-1.81878917E-06 2.81968625E-10-1.63584348E-14    2
-1.68237489E+04-3.20700633E+01 1.93823075E+00 3.01465730E-02-2.61053152E-05    3
 1.09463562E-08-1.78312692E-12-1.38166625E+04 1.85042002E+01                   4
HOCH2O     2/16/99 THERMC   1H   3O   2    0G   300.000  5000.000 1452.000     1
 6.39521515E+00 7.43673043E-03-2.50422354E-06 3.84879712E-10-2.21778689E-14    2
-2.41108840E+04-6.63865583E+00 4.11183145E+00 7.53850697E-03 3.77337370E-06    3
-5.38746005E-09 1.45615887E-12-2.28023001E+04 7.46807254E+00                   4
CH3OH             T06/02C   1H  4 O  1    0 G   200.000  6000.00  1000.00      1
 3.52726795E+00 1.03178783E-02-3.62892944E-06 5.77448016E-10-3.42182632E-14    2
-2.60028834E+04 5.16758693E+00 5.65851051E+00-1.62983419E-02 6.91938156E-05    3
-7.58372926E-08 2.80427550E-11-2.56119736E+04-8.97330508E-01-2.41746056E+04    4
CH2OH             IU2/03C  1 H  3 O  1    0 G   200.000  6000.00   1000.00     1
 5.09314370E+00 5.94761260E-03-2.06497460E-06 3.23008173E-10-1.88125902E-14    2
-4.03409640E+03-1.84691493E+00 4.47834367E+00-1.35070310E-03 2.78484980E-05    3
-3.64869060E-08 1.47907450E-11-3.50072890E+03 3.30913500E+00-2.04462770E+03    4
CH3O              IU1/03C  1 H  3 O  1    0 G   200.000  6000.00  1000.00      1
 4.75779238E+00 7.44142474E-03-2.69705176E-06 4.38090504E-10-2.63537098E-14    2
 3.78111940E+02-1.96680028E+00 3.71180502E+00-2.80463306E-03 3.76550971E-05    3
-4.73072089E-08 1.86588420E-11 1.29569760E+03 6.57240864E+00 2.52571660E+03    4
CH3O2H            A 7/05C  1 H  4 O  2    0 G   200.000  6000.00  1000.00      1
 7.76538058E+00 8.61499712E-03-2.98006935E-06 4.68638071E-10-2.75339255E-14    2
-1.82979984E+04-1.43992663E+01 2.90540897E+00 1.74994735E-02 5.28243630E-06    3
-2.52827275E-08 1.34368212E-11-1.68894632E+04 1.13741987E+01-1.52423685E+04    4
CH3O2                   H   3C   1O   2    0G    300.00   5000.00 1000.00      1
 4.80390863E+00 9.95844638E-03-3.85301026E-06 6.84740497E-10-4.58402955E-14    2
-7.47135460E+02 1.45281400E+00 3.62497097E+00 3.59397933E-03 2.26538097E-05    3
-2.95391947E-08 1.11977570E-11 7.93040410E+01 9.96382194E+00                   4
CH2O2H     1/14/ 5 THERMC   1H   3O   2    0G   300.000  5000.000 1357.000     1
 9.10784249E+00 5.27260434E-03-1.88170543E-06 3.00561364E-10-1.77865959E-14    2
 3.77440183E+03-2.11741044E+01 4.47228333E+00 1.33401095E-02-5.92919725E-06    3
 4.44481025E-10 2.12699899E-13 5.67413711E+03 4.72608208E+00                   4
CH4               G 8/99C  1 H  4    0    0 G   200.000  6000.00  1000.00      1
 1.65326226E+00 1.00263099E-02-3.31661238E-06 5.36483138E-10-3.14696758E-14    2
-1.00095936E+04 9.90506283E+00 5.14911468E+00-1.36622009E-02 4.91453921E-05    3
-4.84246767E-08 1.66603441E-11-1.02465983E+04-4.63848842E+00-8.97226656E+03    4
CH3               IU0702C  1 H  3    0    0 G   200.000  6000.00  1000.00      1
 0.29781206E+01 0.57978520E-02-0.19755800E-05 0.30729790E-09-0.17917416E-13    2
 0.16509513E+05 0.47224799E+01 0.36571797E+01 0.21265979E-02 0.54583883E-05    3
-0.66181003E-08 0.24657074E-11 0.16422716E+05 0.16735354E+01 0.17643935E+05    4
CH2               IU3/03C  1 H  2    0    0 G   200.000  6000.00  1000.00      1
 3.14631886E+00 3.03671259E-03-9.96474439E-07 1.50483580E-10-8.57335515E-15    2
 4.60412605E+04 4.72341711E+00 3.71757846E+00 1.27391260E-03 2.17347251E-06    3
-3.48858500E-09 1.65208866E-12 4.58723866E+04 1.75297945E+00 4.70504920E+04    4
CH2(S)            IU6/03C  1 H  2    0    0 G   200.000  6000.00  1000.00      1
 3.13501686E+00 2.89593926E-03-8.16668090E-07 1.13572697E-10-6.36262835E-15    2
 5.05040504E+04 4.06030621E+00 4.19331325E+00-2.33105184E-03 8.15676451E-06    3
-6.62985981E-09 1.93233199E-12 5.03662246E+04-7.46734310E-01 5.15727280E+04    4
CH                IU3/03C  1 H  1    0    0 G   200.000  6000.00  1000.00      1
 0.25209369E+01 0.17653639E-02-0.46147660E-06 0.59289675E-10-0.33474501E-14    2
 0.70946769E+05 0.74051829E+01 0.34897583E+01 0.32432160E-03-0.16899751E-05    3
 0.31628420E-08-0.14061803E-11 0.70612646E+05 0.20842841E+01 0.71658188E+05    4
CH*               073003C   1H   1          G  0300.00   5000.00  1000.00      1
 0.02196223E+02 0.02340381E-01-0.07058201E-05 0.09007582E-09-0.03855040E-13    2
 0.10419559E+06 0.09178373E+02 0.03200202E+02 0.02072875E-01-0.05134431E-04    3
 0.05733890E-07-0.01955533E-10 0.10393714E+06 0.03331587E+02                   4
C                 L 7/88C   1     0    0   0G   200.000  6000.00  1000.00      1
 0.26055830E+01-0.19593434E-03 0.10673722E-06-0.16423940E-10 0.81870580E-15    2
 0.85411742E+05 0.41923868E+01 0.25542395E+01-0.32153772E-03 0.73379223E-06    3
-0.73223487E-09 0.26652144E-12 0.85442681E+05 0.45313085E+01 0.86195097E+05    4
C2H6              G 8/88C   2H 6    0      0G   200.000  6000.00  1000.00      1
 4.04666411E+00 1.53538802E-02-5.47039485E-06 8.77826544E-10-5.23167531E-14    2
-1.24473499E+04-9.68698313E-01 4.29142572E+00-5.50154901E-03 5.99438458E-05    3
-7.08466469E-08 2.68685836E-11-1.15222056E+04 2.66678994E+00-1.00849652E+04    4
C2H5       8/ 4/ 4 THERMC   2H   5    0    0G   300.000  5000.000 1387.000     1
 5.88784390E+00 1.03076793E-02-3.46844396E-06 5.32499257E-10-3.06512651E-14    2
 1.15065499E+04-8.49651771E+00 1.32730217E+00 1.76656753E-02-6.14926558E-06    3
-3.01143466E-10 4.38617775E-13 1.34284028E+04 1.71789216E+01                   4
C2H4              G 1/00C  2 H  4    0    0 G   200.000  6000.00  1000.00      1
 3.99182724E+00 1.04833908E-02-3.71721342E-06 5.94628366E-10-3.53630386E-14    2
 4.26865851E+03-2.69081762E-01 3.95920063E+00-7.57051373E-03 5.70989993E-05    3
-6.91588352E-08 2.69884190E-11 5.08977598E+03 4.09730213E+00 6.31426266E+03    4
C2H3              ATCT/AC  2 H  3    0    0 G   200.000  6000.00  1000.00      1
 4.15026763E+00 7.54021341E-03-2.62997847E-06 4.15974048E-10-2.45407509E-14    2
 3.38566380E+04 1.72812235E+00 3.36377642E+00 2.65765722E-04 2.79620704E-05    3
-3.72986942E-08 1.51590176E-11 3.44749589E+04 7.91510092E+00 3.56701718E+04    4
C2H2              G 1/91C  2 H  2    0    0 G   200.000  6000.00  1000.00      1
 4.65878489E+00 4.88396667E-03-1.60828888E-06 2.46974544E-10-1.38605959E-14    2
 2.57594042E+04-3.99838194E+00 8.08679682E-01 2.33615762E-02-3.55172234E-05    3
 2.80152958E-08-8.50075165E-12 2.64289808E+04 1.39396761E+01 2.74459950E+04    4
C2H               T 5/10C  2 H  1    0    0 G   200.000  6000.00  1000.00      1
 3.66270248E+00 3.82492252E-03-1.36632500E-06 2.13455040E-10-1.23216848E-14    2
 6.71683790E+04 3.92205792E+00 2.89867676E+00 1.32988489E-02-2.80733327E-05    3
 2.89484755E-08-1.07502351E-11 6.70616050E+04 6.18547632E+00 6.83210436E+04    4
CH3CHO            L 8/88C  2 H  4 O   1   0 G   200.000  6000.00  1000.00      1
 0.54041108E+01 0.11723059E-01-0.42263137E-05 0.68372451E-09-0.40984863E-13    2
-0.22593122E+05-0.34807917E+01 0.47294595E+01-0.31932858E-02 0.47534921E-04    3
-0.57458611E-07 0.21931112E-10-0.21572878E+05 0.41030159E+01-0.19987949E+05    4
CH3CO             IU2/03C  2 H  3 O  1    0 G   200.000  6000.00  1000.00      1
 0.53137165E+01 0.91737793E-02-0.33220386E-05 0.53947456E-09-0.32452368E-13    2
-0.36450414E+04-0.16757558E+01 0.40358705E+01 0.87729487E-03 0.30710010E-04    3
-0.39247565E-07 0.15296869E-10-0.26820738E+04 0.78617682E+01-0.12388039E+04    4
CH2CHO            T03/10C  2 H  3 O  1    0 G   200.000  6000.00  1000.00      1
 6.53928338E+00 7.80238629E-03-2.76413612E-06 4.42098906E-10-2.62954290E-14    2
-1.18858659E+03-8.72091393E+00 2.79502600E+00 1.01099472E-02 1.61750645E-05    3
-3.10303145E-08 1.39436139E-11 1.62944975E+02 1.23646657E+01 1.53380440E+03    4
CH2CO                   H   2C   2O   1    0G    300.00   5000.00 1000.00      1
 5.35869367E+00 6.95641586E-03-2.64802637E-06 4.65067592E-10-3.08641820E-14    2
-7.90294013E+03-3.98525731E+00 1.81422511E+00 1.99008590E-02-2.21416008E-05    3
 1.45028521E-08-3.98877068E-12-7.05394926E+03 1.36079359E+01                   4
HCCO              T 4/09H  1 C  2 O  1    0 G   200.000  6000.00  1000.00      1
 5.91479333E+00 3.71408730E-03-1.30137010E-06 2.06473345E-10-1.21476759E-14    2
 1.93596301E+04-5.50567269E+00 1.87607969E+00 2.21205418E-02-3.58869325E-05    3
 3.05402541E-08-1.01281069E-11 2.01633840E+04 1.36968290E+01 2.14444387E+04    4
HCCOH             T12/09C  2 H  2 O  1    0 G   200.000  6000.00  1000.00      1
 6.37509678E+00 5.49429011E-03-1.88136576E-06 2.93803536E-10-1.71771901E-14    2
 8.93277676E+03-8.24498007E+00 2.05541154E+00 2.52003372E-02-3.80821654E-05    3
 3.09890632E-08-9.89799902E-12 9.76872113E+03 1.22271534E+01 1.12217316E+04    4
CH3CO3H    6/26/95 THERMC   2H   4O   3    0G   300.000  5000.000 1391.000     1
 1.25060485E+01 9.47789695E-03-3.30402246E-06 5.19630793E-10-3.04233568E-14    2
-4.59856703E+04-3.79195947E+01 2.24135876E+00 3.37963514E-02-2.53887482E-05    3
 9.67583587E-09-1.49266157E-12-4.24677831E+04 1.70668133E+01                   4
CH3CO3     4/ 3/ 0 THERMC   2H   3O   3    0G   300.000  5000.000 1391.000     1
 1.12522498E+01 8.33652672E-03-2.89014530E-06 4.52781734E-10-2.64354456E-14    2
-2.60238584E+04-2.96370457E+01 3.60373432E+00 2.70080341E-02-2.08293438E-05    3
 8.50541104E-09-1.43846110E-12-2.34205171E+04 1.12014914E+01                   4
CH3CO2     2/14/95 THERMC   2H   3O   2    0G   300.000  5000.000 1395.000     1
 8.54059736E+00 8.32951214E-03-2.84722010E-06 4.41927196E-10-2.56373394E-14    2
-2.97290678E+04-2.03883545E+01 1.37440768E+00 2.49115604E-02-1.74308894E-05    3
 6.24799508E-09-9.09516835E-13-2.72330150E+04 1.81405454E+01                   4
C2H5OH            L 8/88C  2 H  6 O  1    0 G   200.000  6000.00  1000.00      1
 0.65624365E+01 0.15204222E-01-0.53896795E-05 0.86225011E-09-0.51289787E-13    2
-0.31525621E+05-0.94730202E+01 0.48586957E+01-0.37401726E-02 0.69555378E-04    3
-0.88654796E-07 0.35168835E-10-0.29996132E+05 0.48018545E+01-0.28257829E+05    4
PC2H4OH           T12/01C  2 H  5 O  1    0 G   200.000  6000.00  1000.00      1
 7.02824536E+00 1.20037746E-02-4.21306455E-06 6.69471213E-10-3.96371893E-14    2
-5.92493321E+03-9.40355948E+00 4.47893092E+00 7.59782301E-03 2.81794908E-05    3
-4.26953487E-08 1.78878934E-11-4.71446256E+03 6.38921206E+00-2.86833500E+03    4
SC2H4OH           T10/04C  2 H  5 O  1    0 G   200.000  6000.00  1000.00      1
 6.35842302E+00 1.24356276E-02-4.33096839E-06 6.84530381E-10-4.03713238E-14    2
-9.37900432E+03-6.05106112E+00 4.22283250E+00 5.12174798E-03 3.48386522E-05    3
-4.91943637E-08 2.01183723E-11-8.20503939E+03 8.01675700E+00-6.49827831E+03    4
C2H5O             IU2/03C  2 H  5 O  1    0 G   200.000  6000.00  1000.00      1
 0.66889982E+01 0.13125676E-01-0.47038840E-05 0.75858552E-09-0.45413306E-13    2
-0.47457832E+04-0.96983755E+01 0.43074268E+01 0.64147205E-02 0.31139714E-04    3
-0.43314083E-07 0.17276184E-10-0.34027524E+04 0.59025837E+01-0.16357022E+04    4
O2C2H4OH   2/14/95 THERMC   2H   5O   3    0G   300.000  5000.000 1392.000     1
 1.07432659E+01 1.30957787E-02-4.45370088E-06 6.88548738E-10-3.98230113E-14    2
-2.55911274E+04-2.33254953E+01 4.11839445E+00 2.72240632E-02-1.60824430E-05    3
 5.17033408E-09-7.31610168E-13-2.30857785E+04 1.28482112E+01                   4
C2H5O2H    1/14/ 5 THERMC   2H   6O   2    0G   300.000  5000.000 1391.000     1
 1.12305737E+01 1.20482120E-02-3.96730201E-06 6.00754632E-10-3.42657803E-14    2
-2.47977531E+04-3.25607232E+01 1.57329011E+00 3.52379996E-02-2.53203993E-05    3
 9.56802476E-09-1.48167375E-12-2.15278368E+04 1.90472032E+01                   4
C2H5O2            T10/10C  2 H  5 O  2    0 G   200.000  6000.00  1000.00      1
 8.88872432E+00 1.35833179E-02-4.91116949E-06 7.92343362E-10-4.73525704E-14    2
-7.44107388E+03-1.90789836E+01 4.50099327E+00 6.87965342E-03 4.74143971E-05    3
-6.92287127E-08 2.87395324E-11-5.39547911E+03 7.91490068E+00-3.45206633E+03    4
C2H4O2H    1/14/ 5 THERMC   2H   5O   2    0G   300.000  5000.000 1397.000     1
 1.05228954E+01 9.48091381E-03-3.55727763E-06 6.41445994E-10-4.21232247E-14    2
 1.55718322E+03-2.31413632E+01 3.46916874E+00 2.71188626E-02-2.08022550E-05    3
 8.44284845E-09-1.40756215E-12 3.89688270E+03 1.43400726E+01                   4
CH3CHO2H   1/14/ 5 THERMC   2H   5O   2    0G   300.000  5000.000 1385.000     1
 1.06284708E+01 1.01662327E-02-3.34915963E-06 5.07257146E-10-2.89352540E-14    2
-2.15391230E+03-2.60363030E+01 3.91433011E+00 2.52722102E-02-1.62112291E-05    3
 5.45591592E-09-7.57965290E-13 2.38044573E+02 1.02327238E+01                   4
C2H4O1-2          L 8/88C  2 H  4 O  1    0 G   200.000  6000.00  1000.00      1
 0.54887641E+01 0.12046190E-01-0.43336931E-05 0.70028311E-09-0.41949088E-13    2
-0.91804251E+04-0.70799605E+01 0.37590532E+01-0.94412180E-02 0.80309721E-04    3
-0.10080788E-06 0.40039921E-10-0.75608143E+04 0.78497475E+01-0.63304657E+04    4
C2H3O1-2          A 1/05C  2 H  3 O  1    0 G   200.000  6000.00  1000.00      1
 5.60158035E+00 9.17613962E-03-3.28028902E-06 5.27903888E-10-3.15362241E-14    2
 1.71446252E+04-5.47228512E+00 3.58349017E+00-6.02275805E-03 6.32426867E-05    3
-8.18540707E-08 3.30444505E-11 1.85681353E+04 9.59725926E+00 1.97814471E+04    4
CH3COCH3          ATCT AC  3 H  6 O  1    0 G   200.000  6000.00  1000.00      1
 7.29796974E+00 1.75656913E-02-6.31678065E-06 1.02025553E-09-6.10903592E-14    2
-2.95368927E+04-1.27591704E+01 5.55638920E+00-2.83863547E-03 7.05722951E-05    3
-8.78130984E-08 3.40290951E-11-2.78325393E+04 2.31960221E+00-2.58360384E+04    4
CH3COCH2          A10/04C  3 H  5 O  1    0 G   200.000  6000.00  1000.00      1
 7.54410697E+00 1.43443222E-02-5.08381081E-06 8.13200521E-10-4.83673315E-14    2
-7.48672286E+03-1.14792587E+01 4.70187196E+00 5.51653762E-03 4.27505858E-05    3
-5.94680816E-08 2.40685378E-11-5.92845491E+03 7.12932590E+00-4.00985747E+03    4
CH3COCH2O2  2/14/95     C   3H   5O   3    0G   300.000  5000.000 1379.00      1
 1.27690342E+01 1.42554828E-02-4.92821461E-06 7.70448921E-10-4.49110534E-14    2
-2.34798669E+04-3.27155799E+01 5.95535468E+00 2.70255205E-02-1.37385031E-05    3
 3.53735851E-09-4.03922557E-13-2.06679464E+04 5.21436049E+00                   4
CH3COCH2O2H 2/14/95     C   3H   6O   3    0G   300.000  5000.000 1381.00      1
 1.52372810E+01 1.44114651E-02-5.01290009E-06 7.87071229E-10-4.60225784E-14    2
-4.27564444E+04-4.77383784E+01 4.94789761E+00 3.60474432E-02-2.21719933E-05    3
 6.98296874E-09-9.21269260E-13-3.88687178E+04 8.49926130E+00                   4
CH3COCH2O  4/ 3/ 0 THERMC   3H   5O   2    0G   300.000  5000.000 1370.000     1
 1.14637586E+01 1.32124342E-02-4.56580495E-06 7.13897538E-10-4.16281047E-14    2
-2.23833017E+04-3.15127868E+01 3.72927689E+00 2.63943697E-02-1.09796486E-05    3
 8.58185303E-10 3.39474590E-13-1.91551565E+04 1.18505335E+01                   4
C2H3CHO    6/26/95 THERMC   3H   4O   1    0G   300.000  5000.000 1393.000     1
 1.04184959E+01 9.48963321E-03-3.29310529E-06 5.16279203E-10-3.01587291E-14    2
-1.49630281E+04-3.07235061E+01 2.92355162E-01 3.54321417E-02-2.94936324E-05    3
 1.28100124E-08-2.26144108E-12-1.16521584E+04 2.28878280E+01                   4
C2H3CO     4/ 3/ 0 THERMC   3H   3O   1    0G   300.000  5000.000 1402.000     1
 9.37467676E+00 7.91296900E-03-2.67198280E-06 4.11115430E-10-2.36978981E-14    2
 1.92969514E+03-2.40892696E+01 1.36242013E+00 3.15273972E-02-3.00218935E-05    3
 1.48167112E-08-2.87971530E-12 4.25770215E+03 1.72626546E+01                   4
C2H5CHO           T05/10C  3 H  6 O  1    0 G   200.000  6000.00  1000.00      1
 7.44085690E+00 1.77301764E-02-6.34081568E-06 1.02040803E-09-6.09461714E-14    2
-2.60055814E+04-1.44195446E+01 4.24529681E+00 6.68296706E-03 4.93337933E-05    3
-6.71986124E-08 2.67262347E-11-2.41473007E+04 6.90738560E+00-2.22688471E+04    4
C2H5CO            A10/04C  3 H  5 O  1    0 G   200.000  6000.00  1000.00      1
 6.52325448E+00 1.54211952E-02-5.50898157E-06 8.85889862E-10-5.28846399E-14    2
-7.19631634E+03-5.19862218E+00 6.25722402E+00-9.17612184E-03 7.61190493E-05    3
-9.05514997E-08 3.46198215E-11-5.91616484E+03 2.23330599E+00-3.94851891E+03    4
CH2CH2CHO  8/10/ 4 THERMC   3H   5O   1    0G   300.000  5000.000 1363.000     1
 9.96855598E+00 1.61917946E-02-6.64161740E-06 1.15444520E-09-7.21981790E-14    2
-4.16450354E+03-2.73971573E+01 8.36272659E+00-3.90712606E-03 3.59751257E-05    3
-2.69209237E-08 5.98920261E-12-7.55243244E+02-9.53140102E+00                   4
CH3CHCHO   8/10/ 4 THERMC   3H   5O   1    0G   300.000  5000.000 1253.000     1
 8.27772090E+00 1.95687188E-02-8.47575089E-06 1.53249728E-09-9.86441542E-14    2
-8.34456062E+03-2.17652483E+01-2.72811212E+00 3.80354483E-02-1.96782132E-05    3
 5.09554570E-09-7.28789092E-13-3.51122739E+03 4.04496677E+01                   4
CH3OCH3    1/20/11      C   2H   6O   1    0G   300.000  5000.000 1367.000     1
 7.36358679E+00 1.38910153E-02-4.74083257E-06 7.34874498E-10-4.25867578E-14    2
-2.61148074E+04-1.61332876E+01 2.41860337E+00 1.87279640E-02-1.40894592E-06    3
-4.28367822E-09 1.36818123E-12-2.36771735E+04 1.28877967E+01                   4
CH3OCH2    1/20/11      C   2H   5O   1    0G   300.000  5000.000 1389.000     1
 6.73134670E+00 1.18022530E-02-4.00104434E-06 6.17227325E-10-3.56435023E-14    2
-3.34933412E+03-9.40782513E+00 2.19172957E+00 1.90390966E-02-6.81450700E-06    3
 8.63577609E-11 3.23902492E-13-1.38948253E+03 1.62440756E+01                   4
CH3OCH2O2  1/20/11      C   2H   5O   3    0G   300.000  5000.000 1399.000     1
 1.22024149E+01 1.19225104E-02-4.06624713E-06 6.30079576E-10-3.65065312E-14    2
-2.40327175E+04-3.38665462E+01 1.72101041E+00 3.78155492E-02-2.89668870E-05    3
 1.16796117E-08-1.93234479E-12-2.05308597E+04 2.19296296E+01                   4
CH2OCH2O2H 1/20/11      C   2H   5O   3    0G   300.000  5000.000 1419.000     1
 1.51031233E+01 9.18263324E-03-3.15895361E-06 4.92789411E-10-2.87001298E-14    2
-1.96611854E+04-4.85172618E+01 9.08332173E-01 4.47997444E-02-3.69441578E-05    3
 1.48366604E-08-2.32279459E-12-1.50992319E+04 2.66419885E+01                   4
CH3OCH2O2H 1/20/11      C   2H   6O   3    0G   300.000  5000.000 1402.000     1
 1.46617126E+01 1.20544674E-02-4.13604704E-06 6.43721637E-10-3.74188832E-14    2
-4.18896186E+04-4.81293252E+01 7.37369081E-01 4.67410003E-02-3.73051936E-05    3
 1.50735309E-08-2.43781978E-12-3.73260287E+04 2.57932851E+01                   4
CH3OCH2O   2/ 9/96 THERMC   2H   5O   2    0G   300.000  5000.000 2012.000     1
 8.60261845E+00 1.35772195E-02-4.84661602E-06 7.77766193E-10-4.62633624E-14    2
-2.13762444E+04-1.75775023E+01 3.25889339E+00 2.22146359E-02-7.78556340E-06    3
-2.41484158E-10 4.51914496E-13-1.92377212E+04 1.23680069E+01                   4
O2CH2OCH2O2H 1/20/11    C   2H   5O   5    0G   300.000  5000.000 1411.000     1
 1.96207800E+01 9.96131702E-03-3.41480475E-06 5.31364852E-10-3.08902100E-14    2
-3.98679641E+04-6.72721405E+01-1.22579809E-01 6.64376755E-02-6.55340609E-05    3
 3.13441786E-08-5.79042960E-12-3.41530358E+04 3.49112501E+01                   4
HO2CH2OCHO 1/20/11      C   2H   4O   4    0G   300.000  5000.000 1428.000     1
 1.78528337E+01 7.54042388E-03-2.74895624E-06 4.45343367E-10-2.66154007E-14    2
-6.41380252E+04-6.47357373E+01 5.15432996E-01 4.76081860E-02-3.63877925E-05    3
 1.24225089E-08-1.50813145E-12-5.82730214E+04 2.81992694E+01                   4
OCH2OCHO   1/20/11      C   2H   3O   3    0G   300.000  5000.000 1426.000     1
 1.24378042E+01 7.82259106E-03-2.82874305E-06 4.55808935E-10-2.71391601E-14    2
-4.44526361E+04-3.85337353E+01 3.92797655E+00 1.85731220E-02-4.14656828E-07    3
-6.94060480E-09 2.32311215E-12-4.07070844E+04 1.02048630E+01                   4
HOCH2OCO   8/31/99 THERMC   2H   3O   3    0G   300.000  5000.000 1603.000     1
 1.13737391E+01 8.17663898E-03-2.92034021E-06 4.66695616E-10-2.76276823E-14    2
-4.65575743E+04-2.86035265E+01 6.08180801E+00 1.28768359E-02 2.04419418E-06    3
-6.10154921E-09 1.79820559E-12-4.39526183E+04 2.54054449E+00                   4
CH3OCHO           T 6/08C  2 H  4 O  2    0 G   200.000  6000.00  1000.00      1
 6.33360880E+00 1.34851485E-02-4.84305805E-06 7.81719241E-10-4.67917447E-14    2
-4.68316521E+04-6.91542601E+00 5.96757028E+00-9.38085425E-03 7.07648417E-05    3
-8.29932227E-08 3.13522917E-11-4.55713267E+04 7.50341113E-01-4.37330508E+04    4
CH3OCO            T10/07C  2 H  3 O  2    0 G   200.000  6000.00  1000.00      1
 7.00171955E+00 1.01977290E-02-3.65621800E-06 5.89475086E-10-3.52561321E-14    2
-2.26135780E+04-9.05267669E+00 4.75563598E+00 7.80915313E-03 1.62272935E-05    3
-2.41210787E-08 9.42644561E-12-2.15157456E+04 4.78096491E+00-1.96506108E+04    4
CH2OCHO    4/15/ 8 THERMC   2H   3O   2    0G   300.000  5000.000 1442.000     1
 1.00960096E+01 7.19887066E-03-2.59813465E-06 4.18110812E-10-2.48723387E-14    2
-2.36389018E+04-2.71144175E+01 2.31031671E+00 1.80474065E-02-2.71519637E-06    3
-4.60918579E-09 1.70037078E-12-2.02910878E+04 1.71549722E+01                   4
HE                G 5/97HE 1    0    0    0 G   200.000  6000.00  1000.00      1
 2.50000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-7.45375000E+02 9.28723974E-01 2.50000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-7.45375000E+02 9.28723974E-01 0.00000000E+00    4
C3H8              G 2/00C  3 H  8    0    0 G   200.000  6000.00  1000.00      1
 6.66919760E+00 2.06108751E-02-7.36512349E-06 1.18434262E-09-7.06914630E-14    2
-1.62754066E+04-1.31943379E+01 4.21093013E+00 1.70886504E-03 7.06530164E-05    3
-9.20060565E-08 3.64618453E-11-1.43810883E+04 5.61004451E+00-1.25900384E+04    4
NC3H7             A 5/05C  3 H  7    0    0 G   200.000  6000.00  1000.00      1
 6.49636579E+00 1.77337992E-02-6.24898046E-06 9.95389495E-10-5.90199770E-14    2
 8.85973885E+03-8.56389710E+00 4.08211458E+00 5.23240341E-03 5.13554466E-05    3
-6.99343598E-08 2.81819493E-11 1.04074558E+04 8.39534919E+00 1.21859256E+04    4
IC3H7             A 5/05C  3 H  7    0    0 G   200.000  6000.00  1000.00      1
 5.30597255E+00 1.89854588E-02-6.74315384E-06 1.07993730E-09-6.42785036E-14    2
 7.78748910E+03-2.23233935E+00 5.47421257E+00-8.42536682E-03 8.04607759E-05    3
-9.49287824E-08 3.59830971E-11 9.04939013E+03 3.40542323E+00 1.08473019E+04    4
C3H6              G 2/00C  3 H  6    0    0 G   200.000  6000.00  1000.00      1
 6.03870234E+00 1.62963931E-02-5.82130800E-06 9.35936829E-10-5.58603143E-14    2
-7.41715057E+02-8.43825992E+00 3.83464468E+00 3.29078952E-03 5.05228001E-05    3
-6.66251176E-08 2.63707473E-11 7.88717123E+02 7.53408013E+00 2.40543339E+03    4
C3H5-A            PD5/98C   3H   5    0    0G   300.000  5000.000 1404.000     1
 8.71682542E+00 1.08257699E-02-3.63655884E-06 5.57706282E-10-3.20793321E-14    2
 1.64375315E+04-2.39184681E+01-4.35181829E-01 3.40776627E-02-2.66098022E-05    3
 1.09853986E-08-1.85107479E-12 1.94181924E+04 2.45509858E+01                   4
C3H5-T            PD5/98C   3H   5    0    0G   300.000  5000.000 1389.000     1
 8.25977858E+00 1.14281582E-02-3.89051874E-06 6.02061188E-10-3.48497868E-14    2
 2.64682815E+04-1.97010509E+01 1.12339597E+00 2.68562417E-02-1.65102273E-05    3
 5.28890293E-09-7.08002939E-13 2.91053720E+04 1.91241364E+01                   4
C3H5-S            PD5/98C   3H   5    0    0G   300.000  5000.000 1394.000     1
 8.30447254E+00 1.13525433E-02-3.85583517E-06 5.95730442E-10-3.44434061E-14    2
 2.82273490E+04-2.02359952E+01 5.27650639E-01 2.95749512E-02-2.05159708E-05    3
 7.69163477E-09-1.21882509E-12 3.09544881E+04 2.15637313E+01                   4
C3H4-A            L 8/89C  3 H  4    0    0 G   200.000  6000.00  1000.00      1
 0.63168722E+01 0.11133728E-01-0.39629378E-05 0.63564238E-09-0.37875540E-13    2
 0.20117495E+05-0.10995766E+02 0.26130445E+01 0.12122575E-01 0.18539880E-04    3
-0.34525149E-07 0.15335079E-10 0.21541567E+05 0.10226139E+02 0.22962267E+05    4
C3H4-P            T 2/90H  4 C  3    0    0 G   200.000  6000.00  1000.00      1
 0.60252400E+01 0.11336542E-01-0.40223391E-05 0.64376063E-09-0.38299635E-13    2
 0.19620942E+05-0.86043785E+01 0.26803869E+01 0.15799651E-01 0.25070596E-05    3
-0.13657623E-07 0.66154285E-11 0.20802374E+05 0.98769351E+01 0.22302059E+05    4
C3H3              T 7/11C  3 H  3    0    0 G   200.000  6000.00  1000.000     1
 7.14221719E+00 7.61902211E-03-2.67460030E-06 4.24914904E-10-2.51475443E-14    2
 3.95709594E+04-1.25848690E+01 1.35110873E+00 3.27411291E-02-4.73827407E-05    3
 3.76310220E-08-1.18541128E-11 4.07679941E+04 1.52058598E+01 4.22762135E+04    4
C3H2              T12/00C  3 H  2    0    0 G   200.000  6000.00  1000.00      1
 6.67324762E+00 5.57728845E-03-1.99180164E-06 3.20289156E-10-1.91216272E-14    2
 7.57571184E+04-9.72894405E+00 2.43417332E+00 1.73013063E-02-1.18294047E-05    3
 1.02756396E-09 1.62626314E-12 7.69074892E+04 1.21012230E+01 7.83005132E+04    4
C3H5O      7/20/95 THERMC   3H   5O   1    0G   300.000  5000.000 1380.000     1
 1.02551752E+01 1.14983720E-02-3.84645659E-06 5.88910346E-10-3.38557923E-14    2
 6.26560810E+03-2.77655042E+01 1.19822582E+00 3.05579837E-02-1.80630276E-05    3
 4.86150033E-09-4.19854562E-13 9.58217784E+03 2.15566221E+01                   4
C3H6OOH1-3 7/19/ 0 THERMC   3H   7O   2    0G   300.000  5000.000 1384.000     1
 1.46881564E+01 1.49941200E-02-5.24056505E-06 8.25462711E-10-4.83758952E-14    2
-4.77342863E+03-4.77984492E+01 1.88331465E+00 4.40156051E-02-3.07858462E-05    3
 1.13214862E-08-1.75323184E-12-1.68779168E+02 2.14040621E+01                   4
C3H6OOH1-2 7/19/ 0 THERMC   3H   7O   2    0G   300.000  5000.000 1402.000     1
 1.24605763E+01 1.58889526E-02-5.32742106E-06 8.15818791E-10-4.68723250E-14    2
-4.20305196E+03-3.23858947E+01 2.87774562E+00 3.74166999E-02-2.36058063E-05    3
 7.79930860E-09-1.06042562E-12-7.82368119E+02 1.93941340E+01                   4
C3H6OOH2-1 7/19/ 0 THERMC   3H   7O   2    0G   300.000  5000.000 1407.000     1
 1.42163221E+01 1.43382450E-02-4.78004477E-06 7.29133134E-10-4.17761973E-14    2
-5.67381620E+03-4.35770997E+01 2.09193950E+00 4.69220394E-02-3.90280831E-05    3
 1.72381453E-08-3.07968979E-12-1.89377918E+03 2.00178282E+01                   4
C3H6OOH2-2 7/19/ 0 THERMC   3H   7O   2    0G   300.000  5000.000 1407.000     1
 1.42163221E+01 1.43382450E-02-4.78004477E-06 7.29133134E-10-4.17761973E-14    2
-5.67381620E+03-4.35770997E+01 2.09193950E+00 4.69220394E-02-3.90280831E-05    3
 1.72381453E-08-3.07968979E-12-1.89377918E+03 2.00178282E+01                   4
C3H6OOH1-2O2 7/19/ 0 TRMC   3H   7O   4    0G   300.000  5000.000 1386.000     1
 1.91759159E+01 1.59857013E-02-5.61306378E-06 8.86880495E-10-5.20877040E-14    2
-2.64412115E+04-6.77512936E+01 2.65196584E+00 5.74638149E-02-4.72190867E-05    3
 2.05591557E-08-3.68787387E-12-2.08829371E+04 2.01547955E+01                   4
C3H6OOH1-3O2 7/19/ 0 TRMC   3H   7O   4    0G   300.000  5000.000 1382.000     1
 1.85916698E+01 1.65328553E-02-5.81343626E-06 9.19396939E-10-5.40320702E-14    2
-2.39598698E+04-6.42544402E+01 3.14864588E+00 5.33542571E-02-4.08330611E-05    3
 1.67542220E-08-2.89288326E-12-1.85473645E+04 1.86305431E+01                   4
C3H6OOH2-1O2 7/19/ 0 TRMC   3H   7O   4    0G   300.000  5000.000 1386.000     1
 1.91759159E+01 1.59857013E-02-5.61306378E-06 8.86880495E-10-5.20877040E-14    2
-2.64412115E+04-6.77512936E+01 2.65196584E+00 5.74638149E-02-4.72190867E-05    3
 2.05591557E-08-3.68787387E-12-2.08829371E+04 2.01547955E+01                   4
NC3H7O            T07/10C  3 H  7 O  1    0 G   200.000  6000.00  1000.00      1
 8.38041157E+00 1.95206120E-02-6.97374143E-06 1.12144919E-09-6.69467831E-14    2
-8.48625211E+03-1.89916219E+01 4.21934640E+00 7.38556641E-03 6.02825529E-05    3
-8.38680247E-08 3.39623435E-11-6.23491852E+03 8.08139850E+00-4.26576768E+03    4
IC3H7O     8/ 9/ 4 THERMC   3H   7O   1    0G   300.000  5000.000 1393.000     1
 1.23135031E+01 1.38062606E-02-4.91585531E-06 8.21075632E-10-5.07493001E-14    2
-1.24717023E+04-4.17270532E+01-8.18260771E-01 4.68807147E-02-3.74369377E-05    3
 1.55917264E-08-2.64308171E-12-8.15153216E+03 2.79483196E+01                   4
NC3H7O2H          T02/10C  3 H  8 O  2    0 G   200.000  6000.00  1000.00      1
 1.04115631E+01 2.13763889E-02-7.55819870E-06 1.20207180E-09-7.11798090E-14    2
-2.68935445E+04-2.35428789E+01 7.08977756E+00-4.86163264E-03 1.03253531E-04    3
-1.33200956E-07 5.30799252E-11-2.44194556E+04 1.74859215E+00-2.18476548E+04    4
IC3H7O2H   7/19/ 0 THERMC   3H   8O   2    0G   300.000  5000.000 1389.000     1
 1.57046391E+01 1.65924516E-02-5.77250934E-06 9.06453070E-10-5.30084111E-14    2
-3.23268564E+04-5.71735156E+01 5.19265570E-01 5.32111228E-02-4.05156892E-05    3
 1.63346713E-08-2.73751233E-12-2.71048486E+04 2.40815065E+01                   4
NC3H7O2           T04/10C  3 H  7 O  2    0 G   200.000  6000.00  1000.00      1
 9.24489759E+00 2.14800809E-02-7.69335773E-06 1.23945160E-09-7.40911693E-14    2
-9.81187945E+03-2.20401438E+01 6.99488957E+00-7.50355088E-03 1.01250579E-04    3
-1.25012534E-07 4.84675978E-11-7.53004240E+03-2.03740242E+00-5.10764916E+03    4
IC3H7O2    7/19/ 0 THERMC   3H   7O   2    0G   300.000  5000.000 1388.000     1
 1.32493493E+01 1.64082190E-02-5.67432062E-06 8.87336340E-10-5.17361535E-14    2
-1.44109855E+04-4.29066213E+01 1.49941639E+00 4.43081205E-02-3.22414456E-05    3
 1.29687136E-08-2.23370569E-12-1.02587980E+04 2.02336490E+01                   4
C3H6O1-3          A11/04C  3 H  6 O  1    0 G   200.000  6000.00  1000.00      1
 6.80716906E+00 1.88824545E-02-6.79082475E-06 1.09713919E-09-6.57154952E-14    2
-1.36547629E+04-1.35382154E+01 5.15283752E+00-1.86401716E-02 1.29980652E-04    3
-1.58629974E-07 6.20668783E-11-1.13243512E+04 4.73561224E+00-9.75233898E+03    4
C3H6O1-2          A01/05C  3 H  6 O  1    0 G   200.000  6000.00  1000.00      1
 8.01491079E+00 1.73919953E-02-6.26027968E-06 1.01188256E-09-6.06239111E-14    2
-1.51980838E+04-1.88279964E+01 3.42806676E+00 6.25176642E-03 6.13196311E-05    3
-8.60387185E-08 3.51371393E-11-1.28446646E+04 1.04244994E+01-1.11564001E+04    4
C3KET12    7/19/ 0 THERMC   3H   6O   3    0G   300.000  5000.000 1388.000     1
 1.70756225E+01 1.31013491E-02-4.61949408E-06 7.31991329E-10-4.30788679E-14    2
-4.17008637E+04-5.95778952E+01 1.10507238E+00 5.27396706E-02-4.31805774E-05    3
 1.81618292E-08-3.10535568E-12-3.63627536E+04 2.54111636E+01                   4
C3KET13    7/19/ 0 THERMC   3H   6O   3    0G   300.000  5000.000 1379.000     1
 1.58927479E+01 1.40990923E-02-4.96118851E-06 7.84992198E-10-4.61488928E-14    2
-3.93774829E+04-5.26049341E+01 3.55241022E+00 4.18720270E-02-2.94550370E-05    3
 1.09982900E-08-1.75045977E-12-3.48902671E+04 1.42082894E+01                   4
C3KET21    7/19/ 0 THERMC   3H   6O   3    0G   300.000  5000.000 1371.000     1
 1.56377776E+01 1.44059342E-02-5.08808082E-06 8.07076119E-10-4.75295650E-14    2
-4.30657975E+04-5.13105869E+01 4.55686367E+00 3.57076837E-02-1.94712054E-05    3
 4.70695431E-09-3.69753807E-13-3.86710975E+04 9.97761694E+00                   4
C3H51-2A3OOH 8/26/3 THRMC   3H   7O   4    0G   300.000  5000.000 1386.000     1
 2.12378169E+01 1.39519596E-02-4.94539222E-06 7.86381389E-10-4.63925564E-14    2
-1.92864584E+04-7.69636561E+01 2.55619708E+00 6.13504487E-02-5.23205391E-05    3
 2.28208029E-08-4.02231508E-12-1.31353414E+04 2.21043799E+01                   4
C3H52-1A3OOH 8/26/3 THRMC   3H   7O   4    0G   300.000  5000.000 1379.000     1
 2.02817964E+01 1.48155431E-02-5.25503386E-06 8.35963453E-10-4.93308915E-14    2
-1.80085066E+04-7.22688262E+01 4.12253742E+00 5.19553611E-02-3.83733727E-05    3
 1.45851637E-08-2.29820536E-12-1.22759164E+04 1.48367359E+01                   4
C3H6OH     1/ 7/98 THERMC   3H   7O   1    0G   300.000  5000.000 1674.000     1
 9.31287816E+00 1.67579212E-02-5.75555480E-06 9.00584362E-10-5.26566836E-14    2
-1.20169635E+04-1.95011064E+01 1.20494302E+00 3.30857885E-02-1.63893637E-05    3
 3.18103918E-09-6.84229288E-14-9.12961720E+03 2.47155202E+01                   4
HOC3H6O2   1/ 7/98 THERMC   3H   7O   3    0G   300.000  5000.000 1397.000     1
 1.42691004E+01 1.71837825E-02-5.83419536E-06 9.00994191E-10-5.20716210E-14    2
-3.14501750E+04-4.15295035E+01 3.06954289E+00 4.43105640E-02-3.18636260E-05    3
 1.26409287E-08-2.12751901E-12-2.75893676E+04 1.83891218E+01                   4
CH3CHCO   03/03/95 THERMC   3H   4O   1    0G   300.000  5000.000 1400.00      1
 1.00219123E+01 9.56966300E-03-3.26221644E-06 5.05231706E-10-2.92593257E-14    2
-1.42482738E+04-2.77829973E+01 1.48380119E+00 3.22203013E-02-2.70250033E-05    3
 1.20499164E-08-2.18365931E-12-1.15276540E+04 1.71552068E+01                   4
AC3H5OOH   7/20/98 THERMC   3H   6O   2    0G   300.000  5000.000 1394.000     1
 1.36837693E+01 1.33968049E-02-4.61533631E-06 7.19988958E-10-4.19109988E-14    2
-1.33165248E+04-4.31904193E+01 2.43934647E+00 4.02070638E-02-2.95322679E-05    3
 1.14715600E-08-1.85170511E-12-9.43679906E+03 1.70549969E+01                   4
C2H3OOH    4/18/ 8 THERMC   2H   4O   2    0G   300.000  5000.000 1397.000     1
 1.15749951E+01 8.09909174E-03-2.81808668E-06 4.42697954E-10-2.58998042E-14    2
-8.84852664E+03-3.43859117E+01 1.35644398E+00 3.37002447E-02-2.75988500E-05    3
 1.14222854E-08-1.89488886E-12-5.49996692E+03 1.98354466E+01                   4
C4H10      8/ 4/ 4 THERMC   4H  10    0    0G   300.000  5000.000 1392.000     1
 1.24940183E+01 2.17726258E-02-7.44272215E-06 1.15487023E-09-6.69712949E-14    2
-2.18403437E+04-4.45558921E+01-4.55756824E-01 4.80323389E-02-2.65497552E-05    3
 6.92544700E-09-6.38317504E-13-1.68960904E+04 2.64870966E+01                   4
PC4H9      8/ 4/ 4 THERMC   4H   9    0    0G   300.000  5000.000 1391.000     1
 1.20779744E+01 1.96264778E-02-6.71302199E-06 1.04206424E-09-6.04469282E-14    2
 3.22550473E+03-3.87719384E+01 3.20730933E-01 4.34654454E-02-2.40584970E-05    3
 6.28245308E-09-5.80113166E-13 7.71490893E+03 2.57301085E+01                   4
SC4H9      8/ 4/ 4 THERMC   4H   9    0    0G   300.000  5000.000 1381.000     1
 1.16934304E+01 1.96402287E-02-6.65306517E-06 1.02631895E-09-5.92826294E-14    2
 1.96382429E+03-3.61626672E+01 8.49159986E-01 3.82085320E-02-1.49626797E-05    3
 2.04499211E-10 8.24254437E-13 6.38832956E+03 2.44466606E+01                   4
C4H8-1            T05/09C  4 H  8    0    0 G   200.000  6000.00  1000.00      1
 7.86795262E+00 2.24448843E-02-8.07705438E-06 1.30179988E-09-7.77958472E-14    2
-4.23853340E+03-1.65662549E+01 5.13226136E+00 5.33862838E-03 6.02928960E-05    3
-7.60364685E-08 2.87324693E-11-2.16718358E+03 3.82936810E+00-3.72842176E+00    4
C4H8-2            T 5/09C  4 H  8    0    0 G   200.000  6000.00  1000.00      1
 7.89114667E+00 2.24970532E-02-8.12143779E-06 1.31273568E-09-7.84451632E-14    2
-5.51643171E+03-1.76436027E+01 5.57278967E+00 3.76541017E-03 6.52226708E-05    3
-8.30909522E-08 3.20311342E-11-3.60128327E+03 5.37796708E-01-1.34523863E+03    4
C4H71-1           T05/04C  4 H  7    0    0 G   200.000  6000.00  1000.00      1
 8.15646382E+00 1.90308835E-02-6.73262214E-06 1.07333098E-09-6.36886441E-14    2
 2.55826427E+04-1.61428872E+01 4.19857522E+00 1.19616999E-02 4.23864923E-05    3
-6.30299109E-08 2.59475110E-11 2.75256555E+04 8.57181248E+00 2.95712937E+04    4
C4H71-2           T05/04C  4 H  7    0    0 G   200.000  6000.00  1000.00      1
 8.16688868E+00 1.95680375E-02-6.95694878E-06 1.11504166E-09-6.64079384E-14    2
 2.37537003E+04-1.77041242E+01 3.77145965E+00 1.46544157E-02 3.70080802E-05    3
-5.72714455E-08 2.36641011E-11 2.58014506E+04 9.11906641E+00 2.78022108E+04    4
C4H71-3           T05/04C  4 H  7    0    0 G   200.000  6000.00  1000.00      1
 8.08107449E+00 1.95526544E-02-6.93149115E-06 1.10889183E-09-6.59584410E-14    2
 1.22822959E+04-1.67137903E+01 4.54746808E+00 4.63771460E-03 6.61340221E-05    3
-8.97456502E-08 3.61716165E-11 1.43843217E+04 7.30313471E+00 1.63702936E+04    4
C4H71-4           T05/04C  4 H  7    0    0 G   200.000  6000.00  1000.00      1
 8.49073768E+00 1.91056974E-02-6.74370664E-06 1.07343267E-09-6.36251837E-14    2
 2.04659294E+04-1.74555814E+01 5.07355313E+00 5.27619329E-03 6.23441322E-05    3
-8.54203458E-08 3.45890031E-11 2.24615054E+04 5.60318035E+00 2.46070249E+04    4
C4H72-2           T05/04C  4 H  7    0    0 G   200.000  6000.00  1000.00      1
 7.26612168E+00 1.99858497E-02-7.12030976E-06 1.14276142E-09-6.81206632E-14    2
 2.31915554E+04-1.09941637E+01 7.61389036E+00-9.06922602E-03 8.28486476E-05    3
-9.61203624E-08 3.59333528E-11 2.44971584E+04-5.90519467E+00 2.69231159E+04    4
C4H6              H6W/94C   4H   6    0    0G   300.000  5000.000 1395.000     1
 1.04518247E+01 1.45471475E-02-4.94228994E-06 7.63833067E-10-4.41755383E-14    2
 8.02177132E+03-3.33939064E+01-7.89604392E-01 4.13361127E-02-2.97167286E-05    3
 1.13512399E-08-1.80261184E-12 1.18902568E+04 2.68208195E+01                   4
PC4H9O2H   7/19/ 0 THERMC   4H  10O   2    0G   300.000  5000.000 1387.000     1
 1.82687454E+01 2.16940079E-02-7.54629828E-06 1.18484806E-09-6.92818498E-14    2
-3.39441633E+04-6.84816300E+01 6.34644286E-01 6.20007657E-02-4.34477749E-05    3
 1.61407616E-08-2.53121507E-12-2.76345805E+04 2.67026090E+01                   4
SC4H9O2H   7/19/ 0 THERMC   4H  10O   2    0G   300.000  5000.000 1390.000     1
 1.88587916E+01 2.11200987E-02-7.33205568E-06 1.14969842E-09-6.71656991E-14    2
-3.64236058E+04-7.20026458E+01 3.40587657E-01 6.52078069E-02-4.84840460E-05    3
 1.91011830E-08-3.13833073E-12-3.00007960E+04 2.72835451E+01                   4
PC4H9O2    7/19/ 0 THERMC   4H   9O   2    0G   300.000  5000.000 1385.000     1
 1.57845448E+01 2.15210910E-02-7.44909017E-06 1.16558071E-09-6.79885609E-14    2
-1.60146054E+04-5.40388525E+01 1.94363650E+00 5.15513163E-02-3.28284400E-05    3
 1.13064860E-08-1.70118606E-12-1.08358103E+04 2.13503149E+01                   4
SC4H9O2    7/19/ 0 THERMC   4H   9O   2    0G   300.000  5000.000 1389.000     1
 1.64031135E+01 2.09361006E-02-7.23393011E-06 1.13058996E-09-6.58938667E-14    2
-1.85074517E+04-5.77331636E+01 1.32689044E+00 5.62785583E-02-4.01717786E-05    3
 1.57120967E-08-2.62948443E-12-1.31557057E+04 2.34069659E+01                   4
PC4H9O     8/ 9/ 4 THERMC   4H   9O   1    0G   300.000  5000.000 1403.000     1
 1.49315588E+01 1.95927054E-02-6.66958265E-06 1.03222635E-09-5.97583630E-14    2
-1.46178979E+04-5.25561919E+01-4.99964924E-01 5.37157310E-02-3.44426650E-05    3
 1.08145957E-08-1.29600044E-12-9.11644218E+03 3.09183423E+01                   4
SC4H9O     8/ 9/ 4 THERMC   4H   9O   1    0G   300.000  5000.000 1679.000     1
 1.43323395E+01 2.04542365E-02-7.12271896E-06 1.12545447E-09-6.62697853E-14    2
-1.60006806E+04-5.02030895E+01-4.09000900E-01 5.38573427E-02-3.39105695E-05    3
 1.01023834E-08-1.11268025E-12-1.11109627E+04 2.88554742E+01                   4
C4H7O      4/ 3/ 0 THERMC   4H   7O   1    0G   300.000  5000.000 1395.000     1
 1.53137780E+01 1.43427017E-02-4.81625517E-06 7.39574839E-10-4.26140814E-14    2
-7.29342884E+02-5.52937859E+01-1.60619192E+00 5.58562682E-02-4.35595767E-05    3
 1.70589279E-08-2.65635180E-12 4.85090326E+03 3.47112559E+01                   4
C4H8O1-2   4/ 3/ 0 THERMC   4H   8O   1    0G   300.000  5000.000 1399.000     1
 1.39197290E+01 1.85551492E-02-6.36014179E-06 9.88844645E-10-5.74274779E-14    2
-2.09452548E+04-5.06788231E+01-2.42033073E+00 5.79308508E-02-4.30236499E-05    3
 1.66679793E-08-2.64714350E-12-1.53950880E+04 3.66425242E+01                   4
C4H8O1-3   1/22/95 THERMC   4H   8O   1    0G   300.000  5000.000 1371.000     1
 1.54227092E+01 1.70211052E-02-6.06347951E-06 9.67354762E-10-5.71992419E-14    2
-2.20194174E+04-6.13871862E+01-2.53690104E+00 5.43995707E-02-3.43390305E-05    3
 1.01079922E-08-1.10262736E-12-1.52980680E+04 3.67400719E+01                   4
C4H8O1-4   1/22/95 THERMC   4H   8O   1    0G   300.000  5000.000 1361.000     1
 1.42360731E+01 1.81176105E-02-6.46263809E-06 1.03194372E-09-6.10557331E-14    2
-2.99478670E+04-5.52081041E+01-3.28505561E+00 5.04800902E-02-2.51998984E-05    3
 3.65743744E-09 3.94863161E-13-2.30067422E+04 4.19349253E+01                   4
C4H8O2-3   1/22/95 THERMC   4H   8O   1    0G   300.000  5000.000 1384.000     1
 1.58263859E+01 1.64400938E-02-5.80680311E-06 9.21146000E-10-5.42511002E-14    2
-2.35334573E+04-6.34844562E+01-2.98701197E+00 6.32678880E-02-5.20855777E-05    3
 2.24064364E-08-3.95416618E-12-1.71957196E+04 3.66920390E+01                   4
PC4H8OH    2/12/ 9 THERMC   4H   9O   1    0G   300.000  5000.000 1503.000     1
 1.40357398E+01 1.94173155E-02-6.50230141E-06 9.95481694E-10-5.72034525E-14    2
-1.67631276E+04-4.41162528E+01 1.20329680E+00 4.40218297E-02-2.12295754E-05    3
 3.03714993E-09 3.72027554E-13-1.18622440E+04 2.65515175E+01                   4
SC4H8OH    2/12/ 9 THERMC   4H   9O   1    0G   300.000  5000.000 1392.000     1
 1.48421985E+01 1.78435665E-02-6.16709050E-06 1.00443458E-09-6.10697983E-14    2
-1.81714637E+04-4.96976895E+01-1.04565044E+00 5.72423420E-02-4.43109142E-05    3
 1.80944672E-08-3.02843329E-12-1.28718032E+04 3.48383489E+01                   4
C4H8OH-1O2 6/26/95 THERMC   4H   9O   3    0G   300.000  5000.000 1396.000     1
 1.74383247E+01 2.16778876E-02-7.37772628E-06 1.14128811E-09-6.60391451E-14    2
-3.55892620E+04-5.71247140E+01 2.88497398E+00 5.63287929E-02-3.98403503E-05    3
 1.53891643E-08-2.51940787E-12-3.05246721E+04 2.09293355E+01                   4
C4H8OH-2O2 6/26/95 THERMC   4H   9O   3    0G   300.000  5000.000 1399.000     1
 1.82942871E+01 2.09395389E-02-7.12096934E-06 1.10103094E-09-6.36889768E-14    2
-3.80505855E+04-6.29154326E+01 2.10003504E+00 6.17528218E-02-4.77238541E-05    3
 1.99145784E-08-3.44416275E-12-3.26698755E+04 2.30901271E+01                   4
C4H8OOH1-1 3/27/97 THERMC   4H   9O   2    0G   300.000  5000.000 1379.000     1
 1.80477436E+01 1.92137176E-02-6.66503008E-06 1.04468117E-09-6.10170737E-14    2
-1.23069570E+04-6.33580990E+01 4.36087539E+00 4.46153162E-02-2.14784588E-05    3
 3.14619957E-09 3.03152649E-13-6.89950326E+03 1.24757248E+01                   4
C4H8OOH1-2 7/19/ 0 THERMC   4H   9O   2    0G   300.000  5000.000 1393.000     1
 1.58327906E+01 2.07220436E-02-7.09869028E-06 1.10302045E-09-6.40251984E-14    2
-8.53034314E+03-5.04399828E+01 1.51698234E+00 5.44584331E-02-3.84524319E-05    3
 1.48145523E-08-2.42809434E-12-3.49728423E+03 2.64916926E+01                   4
C4H8OOH1-3 7/19/ 0 THERMC   4H   9O   2    0G   300.000  5000.000 1377.000     1
 1.76442170E+01 1.91706536E-02-6.57168641E-06 1.02246571E-09-5.94304735E-14    2
-1.01859280E+04-6.17115813E+01 1.94106276E+00 5.18789351E-02-3.10411683E-05    3
 8.63568881E-09-8.42841994E-13-4.34315962E+03 2.40230471E+01                   4
C4H8OOH1-4 7/19/ 0 THERMC   4H   9O   2    0G   300.000  5000.000 1386.000     1
 1.78623700E+01 1.95212501E-02-6.80351173E-06 1.06960529E-09-6.26000540E-14    2
-8.87923008E+03-6.34393359E+01 1.45017084E+00 5.72418991E-02-4.06431218E-05    3
 1.52821793E-08-2.42123218E-12-3.02905522E+03 2.50737890E+01                   4
C4H8OOH2-1 7/19/ 0 THERMC   4H   9O   2    0G   300.000  5000.000 1390.000     1
 1.84555673E+01 1.89543719E-02-6.59381457E-06 1.03538370E-09-6.05467101E-14    2
-1.13637100E+04-6.69839138E+01 1.01711681E+00 6.10560866E-02-4.65789185E-05    3
 1.88024138E-08-3.15265575E-12-5.37391474E+03 2.63059691E+01                   4
C4H8OOH2-2 3/27/97 THERMC   4H   9O   2    0G   300.000  5000.000 1383.000     1
 1.63837700E+01 2.04422768E-02-7.04524557E-06 1.09927552E-09-6.39967086E-14    2
-1.45616229E+04-5.33147431E+01 4.40329034E+00 4.30478989E-02-2.14076129E-05    3
 4.28267268E-09-1.27804885E-13-9.79432029E+03 1.30514046E+01                   4
C4H8OOH2-3 7/19/ 0 THERMC   4H   9O   2    0G   300.000  5000.000 1387.000     1
 1.79338472E+01 1.92153623E-02-6.64486961E-06 1.03940007E-09-6.06239862E-14    2
-1.25767913E+04-6.36194089E+01 1.45436266E+00 5.63121286E-02-3.84161425E-05    3
 1.34229297E-08-1.92382914E-12-6.68916116E+03 2.54247554E+01                   4
C4H8OOH2-4 7/19/ 0 THERMC   4H   9O   2    0G   300.000  5000.000 1390.000     1
 1.84555673E+01 1.89543719E-02-6.59381457E-06 1.03538370E-09-6.05467101E-14    2
-1.13637100E+04-6.69839138E+01 1.01711681E+00 6.10560866E-02-4.65789185E-05    3
 1.88024138E-08-3.15265575E-12-5.37391474E+03 2.63059691E+01                   4
C4H8OOH1-2O2 7/19/ 0 TRMC   4H   9O   4    0G   300.000  5000.000 1387.000     1
 2.23244015E+01 2.05474775E-02-7.19076348E-06 1.13361536E-09-6.64744383E-14    2
-3.05468277E+04-8.32666070E+01 2.22400728E+00 7.04994620E-02-5.66978827E-05    3
 2.42627751E-08-4.29715459E-12-2.37391490E+04 2.38371533E+01                   4
C4H8OOH1-3O2 7/19/ 0 TRMC   4H   9O   4    0G   300.000  5000.000 1387.000     1
 2.23244015E+01 2.05474775E-02-7.19076348E-06 1.13361536E-09-6.64744383E-14    2
-3.05468277E+04-8.32666070E+01 2.22400728E+00 7.04994620E-02-5.66978827E-05    3
 2.42627751E-08-4.29715459E-12-2.37391490E+04 2.38371533E+01                   4
C4H8OOH1-4O2 7/19/ 0 TRMC   4H   9O   4    0G   300.000  5000.000 1383.000     1
 2.17116470E+01 2.11216172E-02-7.40101448E-06 1.16772959E-09-6.85139846E-14    2
-2.80483124E+04-7.95885249E+01 3.12351717E+00 6.46725908E-02-4.78357914E-05    3
 1.89656817E-08-3.18025828E-12-2.14664300E+04 2.04322494E+01                   4
C4H8OOH2-1O2 7/19/ 0 TRMC   4H   9O   4    0G   300.000  5000.000 1387.000     1
 2.23244015E+01 2.05474775E-02-7.19076348E-06 1.13361536E-09-6.64744383E-14    2
-3.05468277E+04-8.32666070E+01 2.22400728E+00 7.04994620E-02-5.66978827E-05    3
 2.42627751E-08-4.29715459E-12-2.37391490E+04 2.38371533E+01                   4
C4H8OOH2-3O2 7/19/ 0 TRMC   4H   9O   4    0G   300.000  5000.000 1389.000     1
 2.29951044E+01 1.99238919E-02-6.96326765E-06 1.09677832E-09-6.42747281E-14    2
-3.30095408E+04-8.71461958E+01 2.19248006E+00 7.36763430E-02-6.24428300E-05    3
 2.79371307E-08-5.10126013E-12-2.61773538E+04 2.29568752E+01                   4
C4H8OOH2-4O2 7/19/ 0 TRMC   4H   9O   4    0G   300.000  5000.000 1387.000     1
 2.23244015E+01 2.05474775E-02-7.19076348E-06 1.13361536E-09-6.64744383E-14    2
-3.05468277E+04-8.32666070E+01 2.22400728E+00 7.04994620E-02-5.66978827E-05    3
 2.42627751E-08-4.29715459E-12-2.37391490E+04 2.38371533E+01                   4
NC4KET12   7/19/ 0 THERMC   4H   8O   3    0G   300.000  5000.000 1388.000     1
 2.02458485E+01 1.76440360E-02-6.19054598E-06 9.77688024E-10-5.74053258E-14    2
-4.58141511E+04-7.52145443E+01 8.05387149E-01 6.52375119E-02-5.18373651E-05    3
 2.13454896E-08-3.59860255E-12-3.92395961E+04 2.84908472E+01                   4
NC4KET13   7/19/ 0 THERMC   4H   8O   3    0G   300.000  5000.000 1386.000     1
 1.96430808E+01 1.80940566E-02-6.33063232E-06 9.97860399E-10-5.85076458E-14    2
-4.59588851E+04-7.16905094E+01 2.74883461E+00 5.86936745E-02-4.49605895E-05    3
 1.83200130E-08-3.11765369E-12-4.01065878E+04 1.88072090E+01                   4
NC4KET14   7/19/ 0 THERMC   4H   8O   3    0G   300.000  5000.000 1382.000     1
 1.90283822E+01 1.86604765E-02-6.53616227E-06 1.03102482E-09-6.04833256E-14    2
-4.34678787E+04-6.80210373E+01 3.40797147E+00 5.37386096E-02-3.72613233E-05    3
 1.36862855E-08-2.13798779E-12-3.77919233E+04 1.65580190E+01                   4
NC4KET21   7/19/ 0 THERMC   4H   8O   3    0G   300.000  5000.000 1376.000     1
 1.86231473E+01 1.90969401E-02-6.70745998E-06 1.05994690E-09-6.22564248E-14    2
-4.71929933E+04-6.55477892E+01 4.69785973E+00 4.83859623E-02-3.05576939E-05    3
 1.02705744E-08-1.51713483E-12-4.18665528E+04 1.06715264E+01                   4
NC4KET23   7/19/ 0 THERMC   4H   8O   3    0G   300.000  5000.000 1387.000     1
 1.99512969E+01 1.79558596E-02-6.31230878E-06 9.98217386E-10-5.86636973E-14    2
-4.95585495E+04-7.43071328E+01 4.50575961E-01 6.48862527E-02-5.04446464E-05    3
 2.03085220E-08-3.35952497E-12-4.28779359E+04 3.00153676E+01                   4
NC4KET24   7/19/ 0 THERMC   4H   8O   3    0G   300.000  5000.000 1380.000     1
 1.87707201E+01 1.89490823E-02-6.65182145E-06 1.05080860E-09-6.17069393E-14    2
-4.72319802E+04-6.73335107E+01 2.93007283E+00 5.39296076E-02-3.66164919E-05    3
 1.30880106E-08-1.99245456E-12-4.14118815E+04 1.86567511E+01                   4
C2H5COCH3         T09/10C  4 H  8 O  1    0 G   200.000  6000.000 1000.00      1
 9.29655016E+00 2.29172746E-02-8.22048591E-06 1.32404838E-09-7.91751980E-14    2
-3.34442311E+04-2.04993263E+01 6.61978185E+00 8.51847835E-03 5.10322077E-05    3
-6.58433042E-08 2.49110484E-11-3.15251691E+04-1.09485469E+00-2.88403536E+04    4
C2H5COCH2  4/ 3/ 0 THERMC   4H   7O   1    0G   300.000  5000.000 1383.000     1
 1.42098738E+01 1.57866459E-02-5.50529183E-06 8.65870540E-10-5.06913329E-14    2
-1.41284951E+04-4.87132911E+01 1.54013856E+00 4.39486258E-02-2.97002421E-05    3
 1.05495313E-08-1.58598769E-12-9.50796505E+03 1.99706641E+01                   4
CH2CH2COCH3 6/21/95 THERC   4H   7O   1    0G   300.000  5000.000 1380.00      1
 1.24694368E+01 1.71022143E-02-5.92156726E-06 9.26816806E-10-5.40730504E-14    2
-1.01378242E+04-3.62186375E+01 2.40255609E+00 3.67294268E-02-1.97316510E-05    3
 5.07323216E-09-4.99655275E-13-6.15006886E+03 1.93993386E+01                   4
CH3CHCOCH3 4/ 3/ 0 THERMC   4H   7O   1    0G   300.000  5000.000 1384.000     1
 1.31388032E+01 1.66091073E-02-5.76924215E-06 9.04978165E-10-5.28826527E-14    2
-1.51162098E+04-4.38876580E+01 8.12941079E-01 4.29256944E-02-2.69230252E-05    3
 8.59326807E-09-1.13188129E-12-1.05247481E+04 2.32952685E+01                   4
C2H3COCH3  6/19/95 THERMC   4H   6O   1    0G   300.000  5000.000 1386.00      1
 1.25571995E+01 1.49672645E-02-5.20015351E-06 8.15864365E-10-4.76824406E-14    2
-2.14622958E+04-4.01434299E+01 2.45578501E-01 4.26432049E-02-2.91126822E-05    3
 1.03478392E-08-1.53551381E-12-1.70305379E+04 2.64430799E+01                   4
CH3CHOOCOCH3 6/27/95    C   4H   7O   3    0G   300.000  5000.000 1393.00      1
 1.72170832E+01 1.76740453E-02-6.10387321E-06 9.53711693E-10-5.55757409E-14    2
-3.05280370E+04-5.67959657E+01 1.59405312E+00 5.74729487E-02-4.65071459E-05    3
 2.01816805E-08-3.61175600E-12-2.53445178E+04 2.60857480E+01                   4
CH2CHOOHCOCH3 6/27/95   C   4H   7O   3    0G   300.000  5000.000 1394.00      1
 1.93158016E+01 1.56592602E-02-5.45395604E-06 8.57160086E-10-5.01582885E-14    2
-2.47752201E+04-6.70296581E+01 1.55204769E+00 6.08201262E-02-5.04704383E-05    3
 2.16347587E-08-3.75674081E-12-1.89563540E+04 2.71011896E+01                   4
NC3H7CHO          T05/09 C  4H   8O   1    0G   200.000  6000.000 1000.00      1
 1.02351219E+01 2.32201057E-02-8.46144199E-06 1.37589764E-09-8.27046434E-14    2
-3.00345804E+04-2.82583105E+01 5.30068149E+00 5.00213349E-03 8.12219686E-05    3
-1.07815910E-07 4.25781054E-11-2.71198341E+04 4.93592991E+00-2.47924787E+04    4
NC3H7CO    9/27/95 THERMC   4H   7O   1    0G   300.000  5000.000 1380.00      1
 1.30026331E+01 1.63104877E-02-5.57642899E-06 8.65670629E-10-5.02255667E-14    2
-1.25523385E+04-4.02608515E+01 2.67256826E+00 3.71198825E-02-2.06862859E-05    3
 5.48873888E-09-5.35864183E-13-8.58050888E+03 1.64848950E+01                   4
C3H6CHO-1  9/27/95 THERMC   4H   7O   1    0G   300.000  5000.000 1379.000     1
 1.30322954E+01 1.62418373E-02-5.54388124E-06 8.59723685E-10-4.98459726E-14    2
-6.45915975E+03-3.92399021E+01 2.67672303E+00 3.73064128E-02-2.11281405E-05    3
 5.80472681E-09-6.09688236E-13-2.49714183E+03 1.75750933E+01                   4
C3H6CHO-2 11/15/95 THERMC   4H   7O   1    0G   300.000  5000.000 1682.000     1
 1.11942816E+01 1.81806772E-02-6.35916662E-06 1.00727333E-09-5.93943618E-14    2
-6.86826460E+03-2.80298956E+01 2.95067531E+00 3.34223079E-02-1.45356815E-05    3
 1.67282048E-09 2.62011555E-13-3.79034324E+03 1.74324072E+01                   4
C3H6CHO-3 11/15/95 THERMC   4H   7O   1    0G   300.000  5000.000 1387.000     1
 1.34301738E+01 1.62250792E-02-5.60631713E-06 8.76356273E-10-5.10864241E-14    2
-1.13561098E+04-4.47371262E+01 1.35168659E+00 4.23714083E-02-2.69123192E-05    3
 8.70132567E-09-1.15287455E-12-6.91166610E+03 2.09381509E+01                   4
C2H5CHCO   9/27/95 THERMC   4H   6O   1    0G   300.000  5000.000 1400.00      1
 1.34100537E+01 1.38766678E-02-4.74130143E-06 7.35504188E-10-4.26457752E-14    2
-1.83790837E+04-4.45295352E+01 2.76600655E-01 4.82966593E-02-4.02376928E-05    3
 1.76564254E-08-3.14365357E-12-1.41717351E+04 2.47118671E+01                   4
SC3H5CHO   11/15/95 THERC   4H   6O   1    0G   300.000  5000.000 1390.000     1
 1.31695904E+01 1.42484434E-02-4.90843998E-06 7.65789041E-10-4.45834896E-14    2
-2.04032613E+04-4.43673205E+01 4.35795171E-01 4.48719314E-02-3.36582931E-05    3
 1.33066870E-08-2.17839128E-12-1.60394651E+04 2.37597452E+01                   4
SC3H5CO   11/15/95 THERMC   4H   5O   1    0G   300.000  5000.000 1392.000     1
 1.25514754E+01 1.22521948E-02-4.22382101E-06 6.59184896E-10-3.83818826E-14    2
-4.25349795E+03-4.02864145E+01 1.74191343E+00 3.97229536E-02-3.20061901E-05    3
 1.38227925E-08-2.46272017E-12-6.64428100E+02 1.70762023E+01                   4
IC4H10            G 8/00C  4 H 10    0    0 G   200.000  6000.00  1000.00      1
 9.76991697E+00 2.54997141E-02-9.14142587E-06 1.47328201E-09-8.80799697E-14    2
-2.14052667E+04-3.00329670E+01 4.45479140E+00 8.26058864E-03 8.29886433E-05    3
-1.14647616E-07 4.64569994E-11-1.84593929E+04 4.92740653E+00-1.62354727E+04    4
IC4H9             T 6/04C  4 H  9    0    0 G   200.000  6000.00  1000.00      1
 9.61250942E+00 2.28581786E-02-8.06391309E-06 1.28556553E-09-7.62730799E-14    2
 4.15218608E+03-2.66485099E+01 3.34476784E+00 2.31869650E-02 3.28261040E-05    3
-5.96398514E-08 2.58980820E-11 6.66201200E+03 9.68860372E+00 8.87422590E+03    4
TC4H9             T 6/04C  4 H  9    0    0 G   200.000  6000.00  1000.00      1
 6.72557390E+00 2.53649194E-02-9.05306262E-06 1.45474620E-09-8.67934112E-14    2
 2.57430692E+03-8.89920414E+00 6.45910754E+00-1.02015930E-02 1.06310577E-04    3
-1.25717030E-07 4.75543216E-11 4.43420391E+03 1.30648608E+00 6.61981524E+03    4
IC4H8             T05/09C  4 H  8    0    0 G   200.000  6000.00  1000.00      1
 8.94232121E+00 2.12900129E-02-7.61851464E-06 1.22641473E-09-7.32634442E-14    2
-6.67292929E+03-2.46775148E+01 3.30612340E+00 1.33377057E-02 5.65726066E-05    3
-8.46898088E-08 3.52403438E-11-4.04128388E+03 9.92304633E+00-2.11365432E+03    4
IC4H7             T05/04C  4 H  7    0    0 G   200.000  6000.00  1000.00      1
 8.34970451E+00 1.92508033E-02-6.81360221E-06 1.08484853E-09-6.42422082E-14    2
 1.24406647E+04-1.87060633E+01 2.38739541E+00 2.06784631E-02 2.89299685E-05    3
-5.37553477E-08 2.35670326E-11 1.47584145E+04 1.55529104E+01 1.65497991E+04    4
IC4H9O2    7/19/ 0 THERMC   4H   9O   2    0G   300.000  5000.000 1387.000     1
 1.59741221E+01 2.13534740E-02-7.39001105E-06 1.15624411E-09-6.74408046E-14    2
-1.72329304E+04-5.65302409E+01 1.21434293E+00 5.45388311E-02-3.67001593E-05    3
 1.34131042E-08-2.11741793E-12-1.18482450E+04 2.34153048E+01                   4
TC4H9O2           T04/08C  4 H  9 O  2    0 G   200.000  6000.00  1000.00      1
 1.34566146E+01 2.40864396E-02-8.56308159E-06 1.36853372E-09-8.12706683E-14    2
-1.89690450E+04-4.18792381E+01 4.45494881E+00 2.89185105E-02 3.68274347E-05    3
-7.18116292E-08 3.18779709E-11-1.56103943E+04 9.17831465E+00-1.27983095E+04    4
TC4H8O2H-I 7/19/ 0 THERMC   4H   9O   2    0G   300.000  5000.000 1405.000     1
 1.78060253E+01 1.84952716E-02-6.21268423E-06 9.52753962E-10-5.48010330E-14    2
-1.17555816E+04-6.40180236E+01 1.57469723E+00 6.04648659E-02-4.84991814E-05    3
 2.05236181E-08-3.52974722E-12-6.54190901E+03 2.16852700E+01                   4
IC4H8O2H-I 7/19/ 0 THERMC   4H   9O   2    0G   300.000  5000.000 1388.000     1
 1.80246456E+01 1.93668264E-02-6.74676496E-06 1.06040129E-09-6.20506445E-14    2
-1.00858977E+04-6.57629693E+01 9.94784793E-01 5.89212240E-02-4.25202225E-05    3
 1.61370574E-08-2.55904902E-12-4.08029057E+03 2.58950880E+01                   4
IC4H8O2H-T 7/19/ 0 THERMC   4H   9O   2    0G   300.000  5000.000 1397.000     1
 1.52395012E+01 2.06496983E-02-6.94791927E-06 1.06651097E-09-6.13782754E-14    2
-1.02271199E+04-4.70908585E+01 3.77633001E+00 4.50889269E-02-2.62423875E-05    3
 7.74736900E-09-9.11520393E-13-5.98295842E+03 1.53503399E+01                   4
IC4H8O     7/19/95 THERMC   4H   8O   1    0G   300.000  5000.000 1399.000     1
 1.44624830E+01 1.80562860E-02-6.18008791E-06 9.59941341E-10-5.57132297E-14    2
-2.30230616E+04-5.61190165E+01-2.97373741E+00 6.24618637E-02-5.04348211E-05    3
 2.13345360E-08-3.67382824E-12-1.73274318E+04 3.62336362E+01                   4
CC4H8O     6/29/95 THERMC   4H   8O   1    0G   300.000  5000.000 1401.000     1
 1.35131704E+01 1.91666441E-02-6.53902359E-06 1.01366570E-09-5.87546671E-14    2
-2.00311488E+04-5.22146967E+01-5.27768230E+00 6.52482242E-02-5.00209030E-05    3
 1.97452179E-08-3.15605813E-12-1.37706522E+04 4.78500688E+01                   4
TC4H9O            T08/04C  4 H  9 O  1    0 G   200.000  6000.00  1000.00      1
 1.27371509E+01 2.33707342E-02-8.50516678E-06 1.38519973E-09-8.34398061E-14    2
-1.66940150E+04-4.53156321E+01 2.77057100E+00 2.68033175E-02 4.12718360E-05    3
-7.22054739E-08 3.02642276E-11-1.27079262E+04 1.21532856E+01-1.04543262E+04    4
IC4H9O            A08/04C  4 H  9 O  1    0 G   200.000  6000.00  1000.00      1
 1.16309708E+01 2.47981574E-02-9.01550536E-06 1.46714720E-09-8.83214518E-14    2
-1.37854612E+04-3.81956151E+01 3.80297372E+00 1.56874209E-02 6.81105412E-05    3
-9.83346774E-08 3.95261902E-11-1.00832243E+04 9.78963305E+00-7.82602559E+03    4
IC4H9O2H   7/19/ 0 THERMC   4H  10O   2    0G   300.000  5000.000 1388.000     1
 1.84308794E+01 2.15337606E-02-7.48623965E-06 1.17499240E-09-6.86890788E-14    2
-3.51483277E+04-7.08030846E+01 2.44181899E-01 6.34027841E-02-4.49162379E-05    3
 1.67406877E-08-2.61216478E-12-2.86959808E+04 2.72156229E+01                   4
TC4H9O2H          T02/10C  4 H 10 O  2    0 G   200.000  6000.00  1000.00      1
 1.52702114E+01 2.56462637E-02-9.02796199E-06 1.43759278E-09-8.52381573E-14    2
-3.58539067E+04-5.44966764E+01 3.96033042E+00 4.06267078E-02 1.85652131E-05    3
-5.72128820E-08 2.73014984E-11-3.20467014E+04 7.55565609E+00-2.89963507E+04    4
IC4H7O     4/ 3/ 0 THERMC   4H   7O   1    0G   300.000  5000.000 1386.000     1
 1.33457615E+01 1.61218588E-02-5.44376403E-06 8.38199374E-10-4.83608280E-14    2
 6.11443644E+02-4.36818838E+01 1.74700687E+00 4.07783436E-02-2.44750243E-05    3
 7.06502958E-09-7.51570589E-13 4.86979233E+03 1.94535999E+01                   4
IC4H8OH    2/14/95 THERMC   4H   9O   1    0G   300.000  5000.000 1376.000     1
 1.25605997E+01 2.10637488E-02-7.15019648E-06 1.10439262E-09-6.38428695E-14    2
-1.86203249E+04-3.67889430E+01 3.29612707E+00 3.47649647E-02-1.02505618E-05    3
-2.04641931E-09 1.18879408E-12-1.45627247E+04 1.58606320E+01                   4
IO2C4H8OH  8/23/95 THERMC   4H   9O   3    0G   300.000  5000.000 1395.000     1
 1.79798208E+01 2.13452115E-02-7.29108198E-06 1.13068846E-09-6.55402236E-14    2
-3.85769917E+04-6.23553522E+01 2.88826008E+00 5.80363124E-02-4.26690874E-05    3
 1.71759332E-08-2.91842186E-12-3.33881503E+04 1.83381149E+01                   4
IC3H7CHO   2/22/96 THERMC   4H   8O   1    0G   300.000  5000.000 1391.000     1
 1.37501656E+01 1.83126722E-02-6.28572629E-06 9.78250756E-10-5.68538653E-14    2
-3.26936771E+04-4.77270548E+01-2.73021382E-01 4.89696307E-02-3.12770049E-05    3
 1.00052945E-08-1.27512074E-12-2.76054737E+04 2.83451139E+01                   4
TC3H6CHO   2/22/96 THERMC   4H   7O   1    0G   300.000  5000.000 1389.000     1
 1.31013047E+01 1.66391865E-02-5.68457623E-06 8.81808351E-10-5.11290161E-14    2
-1.30638647E+04-4.42705813E+01 1.87052762E+00 4.14869677E-02-2.66815701E-05    3
 9.01531610E-09-1.27870633E-12-8.97730744E+03 1.66174178E+01                   4
IC3H6CHO   2/22/96 THERMC   4H   7O   1    0G   300.000  5000.000 1390.000     1
 1.33102250E+01 1.62097959E-02-5.57575891E-06 8.69003718E-10-5.05554202E-14    2
-7.62177931E+03-4.25050854E+01 5.21481767E-01 4.43114357E-02-2.86617314E-05    3
 9.30319894E-09-1.20761563E-12-2.99677086E+03 2.68182130E+01                   4
IC3H7CO    2/22/96 THERMC   4H   7O   1    0G   300.000  5000.000 1390.000     1
 1.33305736E+01 1.61873930E-02-5.56711402E-06 8.67575951E-10-5.04696549E-14    2
-1.37307001E+04-4.33958746E+01 5.03452639E-01 4.41607510E-02-2.82139091E-05    3
 8.93548675E-09-1.11327422E-12-9.07755468E+03 2.61991461E+01                   4
TC4H8OOH-IO2 7/19/ 0 TRMC   4H   9O   4    0G   300.000  5000.000 1386.000     1
 2.26382889E+01 2.03246143E-02-7.12390770E-06 1.12425028E-09-6.59732993E-14    2
-3.24406877E+04-8.80387843E+01 2.17782096E+00 7.17785118E-02-5.88836046E-05    3
 2.56759171E-08-4.61678643E-12-2.55622378E+04 2.07846231E+01                   4
IC4H8OOH-IO2 7/19/ 0 TRMC   4H   9O   4    0G   300.000  5000.000 1385.000     1
 2.18969581E+01 2.09637874E-02-7.34664900E-06 1.15926594E-09-6.80225413E-14    2
-2.92664889E+04-8.20540807E+01 2.39424426E+00 6.76572549E-02-5.17083682E-05    3
 2.10796041E-08-3.59960373E-12-2.24787495E+04 2.25029839E+01                   4
IC4H8OOH-TO2 7/19/ 0 TRMC   4H   9O   4    0G   300.000  5000.000 1386.000     1
 2.26382889E+01 2.03246143E-02-7.12390770E-06 1.12425028E-09-6.59732993E-14    2
-3.24406877E+04-8.80387843E+01 2.17782096E+00 7.17785118E-02-5.88836046E-05    3
 2.56759171E-08-4.61678643E-12-2.55622378E+04 2.07846231E+01                   4
IC4KETII   7/19/ 0 THERMC   4H   8O   3    0G   300.000  5000.000 1387.000     1
 1.95143059E+01 1.82377395E-02-6.38908606E-06 1.00801571E-09-5.91440350E-14    2
-4.46884836E+04-7.17167584E+01 1.15501614E+00 6.10622345E-02-4.49711323E-05    3
 1.70514654E-08-2.65948602E-12-3.82747956E+04 2.69612235E+01                   4
IC4KETIT   7/19/ 0 THERMC   4H   8O   3    0G   300.000  5000.000 1388.000     1
 2.09369850E+01 1.71090955E-02-6.01892169E-06 9.52353863E-10-5.59926176E-14    2
-4.77819819E+04-8.27717611E+01 1.14243741E+00 6.33840797E-02-4.73084738E-05    3
 1.77145373E-08-2.67265475E-12-4.09366796E+04 2.34844867E+01                   4
IC4H7OH    4/ 8/97 THERMC   4H   8O   1    0G   300.000  5000.000 1384.000     1
 1.35043419E+01 1.78646968E-02-5.99304371E-06 9.18717641E-10-5.28435302E-14    2
-2.58255688E+04-4.44645715E+01 1.69099899E+00 4.27168891E-02-2.49281695E-05    3
 7.00961522E-09-7.23262828E-13-2.14512334E+04 1.99500833E+01                   4
IC4H6OH    8/19/95 THERMC   4H   7O   1    0G   300.000  5000.000 1390.000     1
 1.40310926E+01 1.55317541E-02-5.32754961E-06 8.28785902E-10-4.81545257E-14    2
-7.69378228E+03-4.76555306E+01 8.63371227E-01 4.68711282E-02-3.43580339E-05    3
 1.33031052E-08-2.13914975E-12-3.14948305E+03 2.29075523E+01                   4
IC3H5CHO   7/19/95 THERMC   4H   6O   1    0G   300.000  5000.000 1396.000     1
 1.36203958E+01 1.37917192E-02-4.73370118E-06 7.36655226E-10-4.20097974E-14    2
-2.00025274E+04-4.73184531E+01 6.27183793E-01 4.66780254E-02-3.74430631E-05    3
 1.58330542E-08-2.73952155E-12-1.57203117E+04 2.16034294E+01                   4
IC3H5CO    4/ 3/ 0 THERMC   4H   5O   1    0G   300.000  5000.000 1397.000     1
 1.30667437E+01 1.16704244E-02-3.99106523E-06 6.19498148E-10-3.59348249E-14    2
-3.36519344E+03-4.35803090E+01 1.85097069E+00 4.18855846E-02-3.62553731E-05    3
 1.65690659E-08-3.05850846E-12 1.70381441E+02 1.53014433E+01                   4
TC3H6OCHO  8/25/95 THERMC   4H   7O   2    0G   300.000  5000.000 1394.00      1
 1.70371287E+01 1.54400645E-02-5.28332886E-06 8.21085347E-10-4.76898429E-14    2
-2.75871941E+04-6.37271230E+01 3.70830259E-01 5.38475661E-02-3.82477565E-05    3
 1.32882237E-08-1.79228730E-12-2.18391262E+04 2.58142112E+01                   4
IC3H6CO   03/03/95 THERMC   4H   6O   1    0G   300.000  5000.000 1397.00      1
 1.32548232E+01 1.40142787E-02-4.78910215E-06 7.42924342E-10-4.30737566E-14    2
-2.00529779E+04-4.44810221E+01 2.28039055E+00 4.17016989E-02-3.25089661E-05    3
 1.37243419E-08-2.40573132E-12-1.63939712E+04 1.38187714E+01                   4
IC4H7OOH   7/19/95 THERMC   4H   8O   2    0G   300.000  5000.000 1392.00      1
 1.69234564E+01 1.78396769E-02-6.14273279E-06 9.57895028E-10-5.57438304E-14    2
-2.00040686E+04-5.94746070E+01 2.99117402E+00 5.03349278E-02-3.56280061E-05    3
 1.33952154E-08-2.11053409E-12-1.51095046E+04 1.54537413E+01                   4
TC3H6OHCHO 8/ 1/95 THERMC   4H   8O   2    0G   300.000  5000.000 1396.00      1
 1.70788996E+01 1.74005554E-02-5.93008112E-06 9.18860909E-10-5.32512140E-14    2
-5.38730427E+04-6.38638754E+01 2.10033500E-01 5.63086284E-02-3.95158669E-05    3
 1.37780428E-08-1.89068805E-12-4.80402638E+04 2.67836070E+01                   4
TC3H6OH    8/ 9/ 4 THERMC   3H   7O   1    0G   300.000  5000.000 1392.000     1
 1.12222277E+01 1.36444398E-02-4.51406709E-06 7.10523275E-10-4.22690392E-14    2
-1.75350136E+04-3.18911926E+01 1.09670360E+00 3.80727565E-02-2.75022497E-05    3
 1.07477493E-08-1.74895773E-12-1.40764487E+04 2.22475799E+01                   4
IC3H5OH    8/ 1/95 THERMC   3H   6O   1    0G   300.000  5000.000 1374.00      1
 1.07381025E+01 1.31698194E-02-4.41529622E-06 6.77009837E-10-3.89608901E-14    2
-2.47298321E+04-3.13634050E+01 1.58376391E+00 3.16215366E-02-1.73664942E-05    3
 4.18927663E-09-2.79899620E-13-2.12643496E+04 1.88313766E+01                   4
TC3H6O2CHO 8/ 2/95 THERMC   4H   7O   3    0G   300.000  5000.000 1386.00      1
 1.85534443E+01 1.68774389E-02-5.90752965E-06 9.31518085E-10-5.46345187E-14    2
-2.85447191E+04-6.82486667E+01 2.17883383E+00 5.41595832E-02-3.83435886E-05    3
 1.38308104E-08-2.04190147E-12-2.27394154E+04 2.00751264E+01                   4
TC3H6O2HCO 8/ 2/95 THERMC   4H   7O   3    0G   300.000  5000.000 1387.00      1
 2.06472678E+01 1.48526500E-02-5.25104875E-06 8.33619219E-10-4.91256069E-14    2
-2.88719869E+04-7.95951389E+01 2.03864428E+00 5.80421003E-02-4.32123528E-05    3
 1.58792094E-08-2.32209543E-12-2.24284673E+04 2.03680990E+01                   4
IC3H5O2HCHO 8/2/95 THERMC   4H   7O   3    0G   300.000  5000.000 1387.00      1
 2.06288832E+01 1.48625539E-02-5.25305276E-06 8.33772951E-10-4.91277401E-14    2
-2.27589076E+04-7.82962888E+01 2.05984770E+00 5.82331716E-02-4.37672100E-05    3
 1.63249918E-08-2.43462051E-12-1.63496250E+04 2.13687921E+01                   4
CH2CCH2OH  9/ 8/95 THERMC   3H   5O   1    0G   300.000  5000.000 1372.00      1
 9.70702027E+00 1.13972660E-02-3.77993962E-06 5.75209277E-10-3.29229125E-14    2
 9.13212884E+03-2.25012933E+01 2.88422544E+00 2.42428071E-02-1.14152268E-05    3
 1.71775334E-09 1.42177454E-13 1.17935615E+04 1.52102335E+01                   4
TC4H8CHO   9/ 7/95 THERMC   5H   9O   1    0G   300.000  5000.000 1397.00      1
 1.79663933E+01 1.94207117E-02-6.67409451E-06 1.03969221E-09-6.04702651E-14    2
-1.33368585E+04-6.79819424E+01-9.58078294E-01 6.42003258E-02-4.70776827E-05    3
 1.75737698E-08-2.64896151E-12-6.86582501E+03 3.33781112E+01                   4
O2C4H8CHO  9/ 7/95 THERMC   5H   9O   3    0G   300.000  5000.000 1395.00      1
 2.12629904E+01 2.14072282E-02-7.38342949E-06 1.15281523E-09-6.71508438E-14    2
-3.16854524E+04-7.99828703E+01 1.91847699E+00 6.67245869E-02-4.80871046E-05    3
 1.78588690E-08-2.71163880E-12-2.49837984E+04 2.38577867E+01                   4
O2HC4H8CO  9/ 7/95 THERMC   5H   9O   3    0G   300.000  5000.000 1394.00      1
 2.38219630E+01 1.91411448E-02-6.67919154E-06 1.05127303E-09-6.15876805E-14    2
-3.23093973E+04-9.42580755E+01 1.82607262E+00 6.93466111E-02-4.93125140E-05    3
 1.69848340E-08-2.26117657E-12-2.46578311E+04 2.41167544E+01                   4
C3H5OH            T06/10C  3 H  6 O  1    0 G   200.000  6000.00  1000.00      1
 8.72477114E+00 1.63942712E-02-5.90852993E-06 9.53262253E-10-5.70318010E-14    2
-1.90496618E+04-1.97198674E+01 3.15011905E+00 1.28538274E-02 4.28438434E-05    3
-6.67818707E-08 2.80408237E-11-1.66413668E+04 1.35066359E+01-1.48710589E+04    4
TIC4H7Q2-I 5/ 6/96 THERMC   4H   9O   4    0G   300.000  5000.000 1400.000     1
 2.33848631E+01 1.87070035E-02-6.44021945E-06 1.00428123E-09-5.84468189E-14    2
-2.61180902E+04-8.76610135E+01 4.48426361E+00 6.61225007E-02-5.27349018E-05    3
 2.18215585E-08-3.66788946E-12-1.98906586E+04 1.26719614E+01                   4
IIC4H7Q2-I 7/15/96 THERMC   4H   9O   4    0G   300.000  5000.000 1394.000     1
 2.30500244E+01 1.92149194E-02-6.66622576E-06 1.04495725E-09-6.10370520E-14    2
-2.32086881E+04-8.39949885E+01 4.93055661E+00 6.05819201E-02-4.23665566E-05    3
 1.49122008E-08-2.10978665E-12-1.68415495E+04 1.36228018E+01                   4
IIC4H7Q2-T 7/15/96 THERMC   4H   9O   4    0G   300.000  5000.000 1377.000     1
 2.15070321E+01 2.05359839E-02-7.12383399E-06 1.11655053E-09-6.52112103E-14    2
-2.51117508E+04-7.43379783E+01 8.16274487E+00 4.34463050E-02-1.76972456E-05    3
 4.88790666E-10 9.03915465E-13-1.96501749E+04 2.62067299E-01                   4
IIC4H7Q2-T 7/15/96 THERMC   4H   9O   4    0G   300.000  5000.000 1377.000     1
 1.59247008E+01 2.59703101E-02-8.86821278E-06 1.37514707E-09-7.97105419E-14    2
-2.60824218E+04-6.16997349E+01-1.67881131E+00 6.41231428E-02-3.96458285E-05    3
 1.23445155E-08-1.53325385E-12-1.96474971E+04 3.39348804E+01                   4
C5H11-1    8/ 4/ 4 THERMC   5H  11    0    0G   300.000  5000.000 1396.000     1
 1.54992372E+01 2.38273176E-02-8.13845161E-06 1.26220569E-09-7.31730066E-14    2
-1.00988975E+03-5.58563592E+01-9.94216435E-01 5.99860809E-02-3.78318587E-05    3
 1.21310895E-08-1.57042863E-12 4.97697538E+03 3.35998032E+01                   4
NC5H12     8/ 4/ 4 THERMC   5H  12    0    0G   300.000  5000.000 1396.000     1
 1.59247008E+01 2.59703101E-02-8.86821278E-06 1.37514707E-09-7.97105419E-14    2
-2.60824218E+04-6.16997349E+01-1.67881131E+00 6.41231428E-02-3.96458285E-05    3
 1.23445155E-08-1.53325385E-12-1.96474971E+04 3.39348804E+01                   4
C5H11-2    8/ 4/ 4 THERMC   5H  11    0    0G   300.000  5000.000 1391.000     1
 1.48744992E+01 2.40593799E-02-8.15587903E-06 1.25867109E-09-7.27223868E-14    2
-2.14733945E+03-5.17907576E+01 7.25187788E-01 4.97343569E-02-2.18806076E-05    3
 2.09007834E-09 6.62752863E-13 3.46418370E+03 2.67485348E+01                   4
C5H11-3    8/ 4/ 4 THERMC   5H  11    0    0G   300.000  5000.000 1391.000     1
 1.48744992E+01 2.40593799E-02-8.15587903E-06 1.25867109E-09-7.27223868E-14    2
-2.14733945E+03-5.24802393E+01 7.25187788E-01 4.97343569E-02-2.18806076E-05    3
 2.09007834E-09 6.62752863E-13 3.46418370E+03 2.60590532E+01                   4
C5H10-1    4/ 7/97 THERMC   5H  10    0    0G   300.000  5000.000 1392.000     1
 1.45851539E+01 2.24072471E-02-7.63348025E-06 1.18188966E-09-6.84385139E-14    2
-1.00898205E+04-5.23683936E+01-1.06223481E+00 5.74218294E-02-3.74486890E-05    3
 1.27364989E-08-1.79609789E-12-4.46546666E+03 3.22739790E+01                   4
C5H10-2    4/ 7/97 THERMC   5H  10    0    0G   300.000  5000.000 1389.000     1
 1.41109267E+01 2.28348272E-02-7.78626835E-06 1.20627491E-09-6.98795983E-14    2
-1.14336507E+04-5.01601163E+01-5.41560551E-01 5.39629918E-02-3.23508738E-05    3
 9.77416037E-09-1.18534668E-12-5.98606169E+03 2.97142748E+01                   4
C5H81-3    3/27/97 THERMC   5H   8    0    0G   300.000  5000.000 1396.000     1
 1.45574490E+01 1.80939266E-02-6.21671892E-06 9.67920254E-10-5.62629326E-14    2
 1.22365462E+03-5.43889766E+01-2.32617433E+00 6.38696042E-02-5.57052591E-05    3
 2.58049480E-08-4.83405924E-12 6.55183321E+03 3.42036513E+01                   4
C5H91-3    4/ 7/97 THERMC   5H   9    0    0G   300.000  5000.000 1392.000     1
 1.41860454E+01 2.07128899E-02-7.06960617E-06 1.09607133E-09-6.35322208E-14    2
 7.00496135E+03-5.14501773E+01-1.38013950E+00 5.57608487E-02-3.70143928E-05    3
 1.26883901E-08-1.78538835E-12 1.25589824E+04 3.26441304E+01                   4
C5H91-4    4/ 7/97 THERMC   5H   9    0    0G   300.000  5000.000 1379.000     1
 1.39904314E+01 1.99962562E-02-6.73105937E-06 1.03447598E-09-5.96148983E-14    2
 1.36075123E+04-4.58753046E+01 2.07302224E-01 4.75322572E-02-2.55232300E-05    3
 5.70570808E-09-2.53926602E-13 1.88300100E+04 2.97527890E+01                   4
C5H91-5    4/ 7/97 THERMC   5H   9    0    0G   300.000  5000.000 1392.000     1
 1.41604486E+01 2.02710046E-02-6.90765357E-06 1.06972742E-09-6.19529514E-14    2
 1.49795090E+04-4.72301324E+01-3.00352280E-01 5.29029897E-02-3.50199571E-05    3
 1.21280172E-08-1.74459793E-12 2.01482388E+04 3.08938514E+01                   4
C5H92-4    4/ 7/97 THERMC   5H   9    0    0G   300.000  5000.000 1389.000     1
 1.37128284E+01 2.11391857E-02-7.22186145E-06 1.12036442E-09-6.49675872E-14    2
 5.66079366E+03-4.92475603E+01-8.61323386E-01 5.23106875E-02-3.19282664E-05    3
 9.73236622E-09-1.17585595E-12 1.10386471E+04 3.00928924E+01                   4
C5H92-5    4/ 7/97 THERMC   5H   9    0    0G   300.000  5000.000 1389.000     1
 1.36885460E+01 2.06966684E-02-7.05980383E-06 1.09401634E-09-6.33885833E-14    2
 1.36345574E+04-4.50306538E+01 2.16350550E-01 4.94614176E-02-2.99438792E-05    3
 9.17728978E-09-1.13613754E-12 1.86282306E+04 2.83575279E+01                   4
C5H9O1-3   4/ 7/97 THERMC   5H   9O   1    0G   300.000  5000.000 1393.000     1
 1.86270165E+01 1.85189638E-02-6.21111137E-06 9.52916260E-10-5.48704082E-14    2
-4.97349374E+03-7.09678919E+01-2.22532588E+00 6.97271843E-02-5.42285799E-05    3
 2.13591167E-08-3.36511599E-12 1.91826163E+03 3.99711270E+01                   4
C5H9O2-4   4/ 7/97 THERMC   5H   9O   1    0G   300.000  5000.000 1387.000     1
 1.86104516E+01 1.87100216E-02-6.31627652E-06 9.73434030E-10-5.62316246E-14    2
-6.59575918E+03-7.05163465E+01-1.66449167E+00 6.51525448E-02-4.57159226E-05    3
 1.55903830E-08-2.04144207E-12 4.10326271E+02 3.84890543E+01                   4
C5H11O-1   4/ 7/97 THERMC   5H  11O   1    0G   300.000  5000.000 1391.000     1
 1.73225378E+01 2.48217999E-02-8.48159842E-06 1.31587304E-09-7.63050620E-14    2
-1.83356880E+04-6.37681611E+01-9.02925873E-02 6.34116550E-02-4.09268668E-05    3
 1.36982820E-08-1.89646466E-12-1.20333690E+04 3.05672313E+01                   4
C5H11O-2   4/ 7/97 THERMC   5H  11O   1    0G   300.000  5000.000 1396.000     1
 1.78183150E+01 2.44541516E-02-8.36505611E-06 1.29863054E-09-7.53356869E-14    2
-2.06350810E+04-6.67615213E+01-4.94527725E-01 6.73149844E-02-4.72324734E-05    3
 1.75936532E-08-2.73651943E-12-1.42372243E+04 3.16370708E+01                   4
C5H11O-3   4/ 7/97 THERMC   5H  11O   1    0G   300.000  5000.000 1396.000     1
 1.78183150E+01 2.44541516E-02-8.36505611E-06 1.29863054E-09-7.53356869E-14    2
-2.06350810E+04-6.74510029E+01-4.94527725E-01 6.73149844E-02-4.72324734E-05    3
 1.75936532E-08-2.73651943E-12-1.42372243E+04 3.09475892E+01                   4
C5H11O2H-1 7/19/ 0 THERMC   5H  12O   2    0G   300.000  5000.000 1387.000     1
 2.14180725E+01 2.62251472E-02-9.10691067E-06 1.42824507E-09-8.34473635E-14    2
-3.80401323E+04-8.39746734E+01 4.74596161E-01 7.38808098E-02-5.12216645E-05    3
 1.87797149E-08-2.90291870E-12-3.05323779E+04 2.91362231E+01                   4
C5H11O2H-2 7/19/ 0 THERMC   5H  12O   2    0G   300.000  5000.000 1390.000     1
 2.21712264E+01 2.55540337E-02-8.86857346E-06 1.39034021E-09-8.12122040E-14    2
-4.06027396E+04-8.84830959E+01-2.68431172E-01 7.90975970E-02-5.89751277E-05    3
 2.33029166E-08-3.83794655E-12-3.28329870E+04 3.17836191E+01                   4
C5H11O2H-3 7/19/ 0 THERMC   5H  12O   2    0G   300.000  5000.000 1390.000     1
 2.21712264E+01 2.55540337E-02-8.86857346E-06 1.39034021E-09-8.12122040E-14    2
-4.06027396E+04-8.84830959E+01-2.68431172E-01 7.90975970E-02-5.89751277E-05    3
 2.33029166E-08-3.83794655E-12-3.28329870E+04 3.17836191E+01                   4
C5H11O2-1  7/19/ 0 THERMC   5H  11O   2    0G   300.000  5000.000 1386.000     1
 1.89702536E+01 2.60355552E-02-9.00706834E-06 1.40888868E-09-8.21618381E-14    2
-2.01253683E+04-6.97477616E+01 1.39788038E+00 6.52788893E-02-4.34224032E-05    3
 1.57151743E-08-2.46631324E-12-1.36791222E+04 2.55411824E+01                   4
C5H11O2-2  7/19/ 0 THERMC   5H  11O   2    0G   300.000  5000.000 1389.000     1
 1.96655539E+01 2.53946113E-02-8.77477373E-06 1.37145913E-09-7.99350015E-14    2
-2.26521255E+04-7.38934310E+01 7.10786402E-01 7.03521821E-02-5.11565299E-05    3
 2.03005197E-08-3.42470585E-12-1.59903126E+04 2.79113132E+01                   4
C5H11O2-3  7/19/ 0 THERMC   5H  11O   2    0G   300.000  5000.000 1389.000     1
 1.96655539E+01 2.53946113E-02-8.77477373E-06 1.37145913E-09-7.99350015E-14    2
-2.26521255E+04-7.38934310E+01 7.10786402E-01 7.03521821E-02-5.11565299E-05    3
 2.03005197E-08-3.42470585E-12-1.59903126E+04 2.79113132E+01                   4
C5H10OOH1-2 7/19/ 0 THRMC   5H  11O   2    0G   300.000  5000.000 1379.000     1
 2.09225281E+01 2.34863057E-02-8.03644420E-06 1.24880724E-09-7.25227776E-14    2
-1.43245680E+04-7.79152904E+01 1.66304681E+00 6.42511734E-02-3.94124754E-05    3
 1.15348101E-08-1.25128422E-12-7.22288006E+03 2.70063739E+01                   4
C5H10OOH1-3 7/19/ 0 THRMC   5H  11O   2    0G   300.000  5000.000 1379.000     1
 2.09225281E+01 2.34863057E-02-8.03644420E-06 1.24880724E-09-7.25227776E-14    2
-1.43245680E+04-7.79152904E+01 1.66304681E+00 6.42511734E-02-3.94124754E-05    3
 1.15348101E-08-1.25128422E-12-7.22288006E+03 2.70063739E+01                   4
C5H10OOH1-4 7/19/ 0 THRMC   5H  11O   2    0G   300.000  5000.000 1379.000     1
 2.09225281E+01 2.34863057E-02-8.03644420E-06 1.24880724E-09-7.25227776E-14    2
-1.43245680E+04-7.79152904E+01 1.66304681E+00 6.42511734E-02-3.94124754E-05    3
 1.15348101E-08-1.25128422E-12-7.22288006E+03 2.70063739E+01                   4
C5H10OOH1-5 7/19/ 0 THRMC   5H  11O   2    0G   300.000  5000.000 1387.000     1
 2.10114488E+01 2.40561226E-02-8.36616955E-06 1.31339875E-09-7.67917194E-14    2
-1.29757849E+04-7.89329903E+01 1.26957212E+00 6.92172253E-02-4.85626715E-05    3
 1.80144791E-08-2.81415382E-12-5.92384799E+03 2.76017751E+01                   4
C5H10OOH2-1 7/19/ 0 THRMC   5H  11O   2    0G   300.000  5000.000 1390.000     1
 2.17441074E+01 2.33958311E-02-8.13002591E-06 1.27566943E-09-7.45598238E-14    2
-1.55260698E+04-8.33092449E+01 5.18861756E-01 7.44934918E-02-5.64622871E-05    3
 2.26488673E-08-3.77612026E-12-8.22372586E+03 3.02858118E+01                   4
C5H10OOH2-3 7/19/ 0 THRMC   5H  11O   2    0G   300.000  5000.000 1388.000     1
 2.10899451E+01 2.37168023E-02-8.19006128E-06 1.27986065E-09-7.45974063E-14    2
-1.66702092E+04-7.91383677E+01 1.27092209E+00 6.82958985E-02-4.63421243E-05    3
 1.61403755E-08-2.30884220E-12-9.58339948E+03 2.79668173E+01                   4
C5H10OOH2-4 7/19/ 0 THRMC   5H  11O   2    0G   300.000  5000.000 1388.000     1
 2.10899451E+01 2.37168023E-02-8.19006128E-06 1.27986065E-09-7.45974063E-14    2
-1.66702092E+04-7.91383677E+01 1.27092209E+00 6.82958985E-02-4.63421243E-05    3
 1.61403755E-08-2.30884220E-12-9.58339948E+03 2.79668173E+01                   4
C5H10OOH2-5 7/19/ 0 THRMC   5H  11O   2    0G   300.000  5000.000 1390.000     1
 2.17441074E+01 2.33958311E-02-8.13002591E-06 1.27566943E-09-7.45598238E-14    2
-1.55260698E+04-8.33092449E+01 5.18861756E-01 7.44934918E-02-5.64622871E-05    3
 2.26488673E-08-3.77612026E-12-8.22372586E+03 3.02858118E+01                   4
C5H10OOH3-1 7/19/ 0 THRMC   5H  11O   2    0G   300.000  5000.000 1390.000     1
 2.17441074E+01 2.33958311E-02-8.13002591E-06 1.27566943E-09-7.45598238E-14    2
-1.55260698E+04-8.33092449E+01 5.18861756E-01 7.44934918E-02-5.64622871E-05    3
 2.26488673E-08-3.77612026E-12-8.22372586E+03 3.02858118E+01                   4
C5H10OOH3-2 7/19/ 0 THRMC   5H  11O   2    0G   300.000  5000.000 1388.000     1
 2.10899451E+01 2.37168023E-02-8.19006128E-06 1.27986065E-09-7.45974063E-14    2
-1.66702092E+04-7.91383677E+01 1.27092209E+00 6.82958985E-02-4.63421243E-05    3
 1.61403755E-08-2.30884220E-12-9.58339948E+03 2.79668173E+01                   4
C5H10O1-2  1/22/95 THERMC   5H  10O   1    0G   300.000  5000.000 1382.000     1
 1.83450823E+01 2.15894287E-02-7.59914917E-06 1.20265688E-09-7.07149348E-14    2
-2.52918816E+04-7.38748127E+01-2.50915891E+00 7.02820905E-02-5.23078154E-05    3
 2.05330738E-08-3.37999472E-12-1.79263879E+04 3.83402738E+01                   4
C5H10O1-3  1/22/95 THERMC   5H  10O   1    0G   300.000  5000.000 1370.000     1
 1.85051134E+01 2.17909650E-02-7.74803799E-06 1.23453810E-09-7.29327086E-14    2
-2.62151881E+04-7.74524221E+01-2.70067147E+00 6.51234466E-02-3.97863209E-05    3
 1.12983558E-08-1.18141056E-12-1.81611984E+04 3.87589334E+01                   4
C5H10O1-4  1/22/95 THERMC   5H  10O   1    0G   300.000  5000.000 1371.000     1
 1.77074517E+01 2.24725523E-02-7.98404192E-06 1.27146816E-09-7.50866945E-14    2
-3.63066445E+04-7.27392560E+01-3.94205066E+00 6.68440102E-02-4.09940878E-05    3
 1.17684771E-08-1.26029870E-12-2.80943137E+04 4.58617150E+01                   4
C5H10O1-5  1/22/95 THERMC   5H  10O   1    0G   300.000  5000.000 1457.000     1
 2.13684109E+01 1.97321411E-02-7.12842160E-06 1.14789888E-09-6.83162787E-14    2
-3.89834904E+04-1.00032176E+02-3.02904503E+00 6.01320166E-02-2.12072490E-05    3
-4.91313274E-09 3.07577547E-12-2.91028862E+04 3.64698785E+01                   4
C5H10O2-3  1/22/95 THERMC   5H  10O   1    0G   300.000  5000.000 1385.000     1
 1.89379846E+01 2.10434849E-02-7.40107577E-06 1.17069402E-09-6.88106356E-14    2
-2.76228814E+04-7.74017673E+01-3.03891874E+00 7.46406721E-02-5.91275018E-05    3
 2.46307903E-08-4.24312686E-12-2.01088998E+04 4.00106761E+01                   4
C5H10O2-4  1/22/95 THERMC   5H  10O   1    0G   300.000  5000.000 1376.000     1
 1.91186278E+01 2.12169126E-02-7.53764833E-06 1.20035780E-09-7.08866585E-14    2
-2.85216189E+04-8.03408390E+01-3.50702064E+00 7.13707278E-02-4.99483546E-05    3
 1.76515898E-08-2.56653255E-12-2.03198734E+04 4.22612571E+01                   4
C5H10OOH1-2O2 7/19/ 0 TMC   5H  11O   4    0G   300.000  5000.000 1387.000     1
 2.55478814E+01 2.50385111E-02-8.74243938E-06 1.37611416E-09-8.06073182E-14    2
-3.46345151E+04-9.91022020E+01 2.53072834E+00 8.12167401E-02-6.33054798E-05    3
 2.63900700E-08-4.58739612E-12-2.67337637E+04 2.39105049E+01                   4
C5H10OOH1-3O2 7/19/ 0 TMC   5H  11O   4    0G   300.000  5000.000 1387.000     1
 2.55478814E+01 2.50385111E-02-8.74243938E-06 1.37611416E-09-8.06073182E-14    2
-3.46345151E+04-9.91022020E+01 2.53072834E+00 8.12167401E-02-6.33054798E-05    3
 2.63900700E-08-4.58739612E-12-2.67337637E+04 2.39105049E+01                   4
C5H10OOH1-4O2 7/19/ 0 TMC   5H  11O   4    0G   300.000  5000.000 1387.000     1
 2.55478814E+01 2.50385111E-02-8.74243938E-06 1.37611416E-09-8.06073182E-14    2
-3.46345151E+04-9.91022020E+01 2.53072834E+00 8.12167401E-02-6.33054798E-05    3
 2.63900700E-08-4.58739612E-12-2.67337637E+04 2.39105049E+01                   4
C5H10OOH1-5O2 7/19/ 0 TMC   5H  11O   4    0G   300.000  5000.000 1385.000     1
 2.48666576E+01 2.56688838E-02-8.97169324E-06 1.41315614E-09-8.28158711E-14    2
-3.21479218E+04-9.51211738E+01 2.81997434E+00 7.72690504E-02-5.67282509E-05    3
 2.23236523E-08-3.71501383E-12-2.43447483E+04 2.35135259E+01                   4
C5H10OOH2-1O2 7/19/ 0 TMC   5H  11O   4    0G   300.000  5000.000 1387.000     1
 2.55478814E+01 2.50385111E-02-8.74243938E-06 1.37611416E-09-8.06073182E-14    2
-3.46345151E+04-9.91022020E+01 2.53072834E+00 8.12167401E-02-6.33054798E-05    3
 2.63900700E-08-4.58739612E-12-2.67337637E+04 2.39105049E+01                   4
C5H10OOH2-3O2 7/19/ 0 TMC   5H  11O   4    0G   300.000  5000.000 1389.000     1
 2.62850175E+01 2.43678422E-02-8.50101950E-06 1.33736519E-09-7.83075048E-14    2
-3.71537284E+04-1.03435286E+02 2.08935173E+00 8.57156954E-02-7.04986902E-05    3
 3.07497216E-08-5.51132533E-12-2.90970365E+04 2.50297599E+01                   4
C5H10OOH2-4O2 7/19/ 0 TMC   5H  11O   4    0G   300.000  5000.000 1389.000     1
 2.62850175E+01 2.43678422E-02-8.50101950E-06 1.33736519E-09-7.83075048E-14    2
-3.71537284E+04-1.03435286E+02 2.08935173E+00 8.57156954E-02-7.04986902E-05    3
 3.07497216E-08-5.51132533E-12-2.90970365E+04 2.50297599E+01                   4
C5H10OOH2-5O2 7/19/ 0 TMC   5H  11O   4    0G   300.000  5000.000 1387.000     1
 2.55478814E+01 2.50385111E-02-8.74243938E-06 1.37611416E-09-8.06073182E-14    2
-3.46345151E+04-9.91022020E+01 2.53072834E+00 8.12167401E-02-6.33054798E-05    3
 2.63900700E-08-4.58739612E-12-2.67337637E+04 2.39105049E+01                   4
C5H10OOH3-1O2 7/19/ 0 TMC   5H  11O   4    0G   300.000  5000.000 1387.000     1
 2.55478814E+01 2.50385111E-02-8.74243938E-06 1.37611416E-09-8.06073182E-14    2
-3.46345151E+04-9.91022020E+01 2.53072834E+00 8.12167401E-02-6.33054798E-05    3
 2.63900700E-08-4.58739612E-12-2.67337637E+04 2.39105049E+01                   4
C5H10OOH3-2O2 7/19/ 0 TMC   5H  11O   4    0G   300.000  5000.000 1389.000     1
 2.62850175E+01 2.43678422E-02-8.50101950E-06 1.33736519E-09-7.83075048E-14    2
-3.71537284E+04-1.03435286E+02 2.08935173E+00 8.57156954E-02-7.04986902E-05    3
 3.07497216E-08-5.51132533E-12-2.90970365E+04 2.50297599E+01                   4
NC5KET12   7/19/ 0 THERMC   5H  10O   3    0G   300.000  5000.000 1389.000     1
 2.34427049E+01 2.21540692E-02-7.74817880E-06 1.22107095E-09-7.15883644E-14    2
-4.99350593E+04-9.09970812E+01 5.64845658E-01 7.74889690E-02-6.00818427E-05    3
 2.42432817E-08-4.02329880E-12-4.21262314E+04 3.12910774E+01                   4
NC5KET13   7/19/ 0 THERMC   5H  10O   3    0G   300.000  5000.000 1387.000     1
 2.27897549E+01 2.26387719E-02-7.89832354E-06 1.24260309E-09-7.27609759E-14    2
-5.00526193E+04-8.71676166E+01 2.53945153E+00 7.08645319E-02-5.32266350E-05    3
 2.12906293E-08-3.56676536E-12-4.29988725E+04 2.14543054E+01                   4
NC5KET14   7/19/ 0 THERMC   5H  10O   3    0G   300.000  5000.000 1387.000     1
 2.27897549E+01 2.26387719E-02-7.89832354E-06 1.24260309E-09-7.27609759E-14    2
-5.00526193E+04-8.71676166E+01 2.53945153E+00 7.08645319E-02-5.32266350E-05    3
 2.12906293E-08-3.56676536E-12-4.29988725E+04 2.14543054E+01                   4
NC5KET15   7/19/ 0 THERMC   5H  10O   3    0G   300.000  5000.000 1383.000     1
 2.21776239E+01 2.31939864E-02-8.09797899E-06 1.27464047E-09-7.46625107E-14    2
-4.75611599E+04-8.35091033E+01 3.22565144E+00 6.57620962E-02-4.52752542E-05    3
 1.64810866E-08-2.54467139E-12-4.06876266E+04 1.90851234E+01                   4
NC5KET21   7/19/ 0 THERMC   5H  10O   3    0G   300.000  5000.000 1379.000     1
 2.17534680E+01 2.36666119E-02-8.28610759E-06 1.30663620E-09-7.66324076E-14    2
-5.12815467E+04-8.09340957E+01 4.56687437E+00 6.01978739E-02-3.82935508E-05    3
 1.29220662E-08-1.89791227E-12-4.47703435E+04 1.29580830E+01                   4
NC5KET23   7/19/ 0 THERMC   5H  10O   3    0G   300.000  5000.000 1387.000     1
 2.31409808E+01 2.24801534E-02-7.87662916E-06 1.24282516E-09-7.29252729E-14    2
-5.36784029E+04-9.00538236E+01 1.09304151E-01 7.75997760E-02-5.94124810E-05    3
 2.36744270E-08-3.89094338E-12-4.57495597E+04 3.32799795E+01                   4
NC5KET24   7/19/ 0 THERMC   5H  10O   3    0G   300.000  5000.000 1385.000     1
 2.25126387E+01 2.29495597E-02-8.02286486E-06 1.26389975E-09-7.40777420E-14    2
-5.38122195E+04-8.63788737E+01 2.19333641E+00 7.04050260E-02-5.15856312E-05    3
 2.00741570E-08-3.28568948E-12-4.66368524E+04 2.29520202E+01                   4
NC5KET25   7/19/ 0 THERMC   5H  10O   3    0G   300.000  5000.000 1382.000     1
 2.19099644E+01 2.35018200E-02-8.22261497E-06 1.29606701E-09-7.59914647E-14    2
-5.13242006E+04-8.27708903E+01 2.76270425E+00 6.58724877E-02-4.45144578E-05    3
 1.58213340E-08-2.38800145E-12-4.43093682E+04 2.11180678E+01                   4
NC5KET31   7/19/ 0 THERMC   5H  10O   3    0G   300.000  5000.000 1382.000     1
 2.17723599E+01 2.36116706E-02-8.25813864E-06 1.30129886E-09-7.62813000E-14    2
-5.13543364E+04-8.16385880E+01 3.14481499E+00 6.64310592E-02-4.75232545E-05    3
 1.85573234E-08-3.11995924E-12-4.46228757E+04 1.89760116E+01                   4
NC5KET32   7/19/ 0 THERMC   5H  10O   3    0G   300.000  5000.000 1387.000     1
 2.29536744E+01 2.26192649E-02-7.91922638E-06 1.24883440E-09-7.32467701E-14    2
-5.36792159E+04-8.86117968E+01 7.24497110E-01 7.71622935E-02-6.10369902E-05    3
 2.55909432E-08-4.44696298E-12-4.60989830E+04 3.00522534E+01                   4
C5H10OH-1  1/14/99 THERMC   5H  11O   1    0G   300.000  5000.000 1371.000     1
 1.75642279E+01 2.33577469E-02-7.81503517E-06 1.19674654E-09-6.88114207E-14    2
-2.11605652E+04-6.19821034E+01 9.51873649E-01 5.58286144E-02-2.87750953E-05    3
 5.54684921E-09 1.10578801E-14-1.48168651E+04 2.93877119E+01                   4
C5H10OH-2  1/14/99 THERMC   5H  11O   1    0G   300.000  5000.000 1390.000     1
 1.72742775E+01 2.39409708E-02-8.07388576E-06 1.24188426E-09-7.15926603E-14    2
-2.31054055E+04-6.11106423E+01 4.68530877E-01 6.05595171E-02-3.75900684E-05    3
 1.16488887E-08-1.41506375E-12-1.70158316E+04 3.00652481E+01                   4
O2C5H10OH-1 1/14/99 THRMC   5H  11O   3    0G   300.000  5000.000 1395.000     1
 2.06059936E+01 2.61750874E-02-8.92270421E-06 1.38184638E-09-8.00235870E-14    2
-4.07496333E+04-7.38943495E+01 2.70461132E+00 6.83289096E-02-4.77921008E-05    3
 1.81238720E-08-2.90871344E-12-3.44822614E+04 2.22673007E+01                   4
O2C5H10OH-2 1/14/99 THRMC   5H  11O   3    0G   300.000  5000.000 1398.000     1
 2.15259930E+01 2.54039694E-02-8.65952886E-06 1.34110440E-09-7.76663740E-14    2
-4.32473477E+04-8.00796638E+01 1.89616952E+00 7.37918569E-02-5.55488679E-05    3
 2.24979959E-08-3.79045894E-12-3.66230283E+04 2.45460172E+01                   4
C6H6              G 6/01C   6H   6    0    0G   200.000  6000.000 1000.000     1
 1.10809576E+01 2.07176746E-02-7.52145991E-06 1.22320984E-09-7.36091279E-14    2
 4.30641035E+03-4.00413310E+01 5.04818632E-01 1.85020642E-02 7.38345881E-05    3
-1.18135741E-07 5.07210429E-11 8.55247913E+03 2.16412893E+01 9.96811598E+03    4
C*CCJC*C   3/1/95  Z&B  C   5H   7    0    0G   300.000  5000.000 1388.000     1
 1.40879309E+01 1.62398907E-02-5.64768950E-06 8.86857524E-10-5.18698993E-14    2
 1.76798698E+04-5.13735038E+01-2.94595603E+00 5.68783623E-02-4.31336497E-05    3
 1.68169537E-08-2.67926433E-12 2.35156925E+04 3.98188778E+01                   4
CC3H4             T12/81C   3H   4    0    0G   300.000  5000.00  1000.00      1
 0.66999931E+01 0.10357372E-01-0.34551167E-05 0.50652949E-09-0.26682276E-13    2
 0.30199051E+05-0.13378770E+02-0.24621047E-01 0.23197215E-01-0.18474357E-05    3
-0.15927593E-07 0.86846155E-11 0.32334137E+05 0.22729762E+02 0.3332728 E+05    4
C4H4              H6W/94C   4H   4    0    0G   300.000  3000.00  1000.00      1
 0.66507092E+01 0.16129434E-01-0.71938875E-05 0.14981787E-08-0.11864110E-12    2
 0.31195992E+05-0.97952118E+01-0.19152479E+01 0.52750878E-01-0.71655944E-04    3
 0.55072423E-07-0.17286228E-10 0.32978504E+05 0.31419983E+02                   4
C4H3-I            AB1/93C   4H   3    0    0G   300.000  3000.00  1000.00      1
 0.90978165E+01 0.92207119E-02-0.33878441E-05 0.49160498E-09-0.14529780E-13    2
 0.56600574E+05-0.19802597E+02 0.20830412E+01 0.40834274E-01-0.62159685E-04    3
 0.51679358E-07-0.17029184E-10 0.58005129E+05 0.13617462E+02                   4
C4H612            A 8/83C   4H   6    0    0G   300.     3000.    1000.0       1
  0.1781557E 02 -0.4257502E-02  0.1051185E-04 -0.4473844E-08  0.5848138E-12    2
  0.1267342E 05 -0.6982662E 02  0.1023467E 01  0.3495919E-01 -0.2200905E-04    3
  0.6942272E-08 -0.7879187E-12  0.1811799E 05  0.1975066E 02  0.1950807E+05    4
C6H5              T04/02C   6H   5    0    0G   200.000  6000.000 1000.        1
 1.08444762E+01 1.73212473E-02-6.29233249E-06 1.02369961E-09-6.16216828E-14    2
 3.55598475E+04-3.53735134E+01 2.10306633E-01 2.04745507E-02 5.89743006E-05    3
-1.01534255E-07 4.47105660E-11 3.95468722E+04 2.52910455E+01 4.08610970E+04    4
C4H2              D11/99C   4H   2    0    0G   300.000  3000.000              1
 0.91576328E+01 0.55430518E-02-0.13591604E-05 0.18780075E-10 0.23189536E-13    2
 0.52588039E+05-0.23711460E+02 0.10543978E+01 0.41626960E-01-0.65871784E-04    3
 0.53257075E-07-0.16683162E-10 0.54185211E+05 0.14866591E+02                   4
C4H3-N            H6W/94C   4H   3    0    0G   300.000  3000.00  1000.00      1
 0.54328279E+01 0.16860981E-01-0.94313109E-05 0.25703895E-08-0.27456309E-12    2
 0.61600680E+05-0.15673981E+01-0.31684113E+00 0.46912100E-01-0.68093810E-04    3
 0.53179921E-07-0.16523005E-10 0.62476199E+05 0.24622559E+02                   4
C4H5-N            H6W/94C   4H   5    0    0G   300.000  3000.00  1000.00      1
 0.98501978E+01 0.10779008E-01-0.13672125E-05-0.77200535E-09 0.18366314E-12    2
 0.38840301E+05-0.26001846E+02 0.16305321E+00 0.39830137E-01-0.34000128E-04    3
 0.15147233E-07-0.24665825E-11 0.41429766E+05 0.23536163E+02                   4
C4H5-I            H6W/94C   4H   5    0    0G   300.000  3000.00  1000.00      1
 0.10229092E+02 0.94850138E-02-0.90406445E-07-0.12596100E-08 0.24781468E-12    2
 0.34642812E+05-0.28564529E+02-0.19932900E-01 0.38005672E-01-0.27559450E-04    3
 0.77835551E-08 0.40209383E-12 0.37496223E+05 0.24394241E+02                   4
CH3CHCHCO         T03/97C   4H   5O   1    0G   200.000  6000.000  1000.0      1
 8.90967920E+00 1.34364140E-02-7.62977390E-07-1.69114810E-09 2.95540440E-13    2
 1.48898740E+03-1.79662460E+01-1.08199860E+00 3.64929760E-02-1.52255950E-05    3
-5.62607170E-18 2.16113750E-21 3.56713230E+03 3.27142550E+01 4.73074990E+03    4
CH2CHCHCHO        T03/97C   4H   5O   1    0G   200.000  6000.000  1000.0      1
 8.90967920E+00 1.34364140E-02-7.62977390E-07-1.69114810E-09 2.95540440E-13    2
 1.48898740E+03-1.79662460E+01-1.08199860E+00 3.64929760E-02-1.52255950E-05    3
-5.62607170E-18 2.16113750E-21 3.56713230E+03 3.27142550E+01 4.73074990E+03    4
C4H6O25           T 3/97C   4H   6O   1    0G   200.000  5000.000  1000.0      1
 8.60658242E+00 2.08310051E-02-8.42229481E-06 1.56717640E-09-1.09391202E-13    2
-1.76177415E+04-2.32464750E+01 2.67053463E+00 4.92586420E-03 8.86967406E-05    3
-1.26219194E-07 5.23991321E-11-1.46572472E+04 1.45722395E+01-1.30831522E+04    4
C2H3CHOCH2        A 8/83C   4H   6O   1    0G   300.     3000.     1000.0      1
-4.72093360E+00 3.91413780E-02-6.52872650E-06-7.68209500E-09 2.51473310E-12    2
 1.75352252E+03 5.17190420E+01 7.97985440E-01 3.44034320E-02-1.24598510E-05    3
-5.18062790E-18 1.99359540E-21-6.48927540E+02 2.18896980E+01 1.00654250E+03    4
C4H5-2            H6W/94C   4H   5    0    0G   300.000  3000.00  1000.00      1
 1.45381710E+01-8.56770560E-03 2.35595240E-05-1.36763790E-08 2.44369270E-12    2
 3.32590950E+04-4.53694970E+01 2.96962800E+00 2.44422450E-02-9.12514240E-06    3
-4.24668710E-18 1.63047280E-21 3.55033160E+04 1.20360510E+01 3.73930550E+04    4
C4H6-2            A 8/83C   4H   6    0    0G   300.     3000.     1000.0      1
  9.0338133E+00  8.2124510E-03  7.1753952E-06 -5.8834334E-09  1.0343915E-12    2
  1.4335068E+04 -2.0985762E+01  2.1373338E+00  2.6486229E-02 -9.0568711E-06    3
 -5.5386397E-19  2.1281884E-22  1.5710902E+04  1.3529426E+01  1.7488676E+04    4
C4H6O23           T 3/97C   4H   6O   1    0G   200.000  5000.000  1000.0      1
 8.60658242E+00 2.08310051E-02-8.42229481E-06 1.56717640E-09-1.09391202E-13    2
-1.32392815E+04-2.32464750E+01 2.67053463E+00 4.92586420E-03 8.86967406E-05    3
-1.26219194E-07 5.23991321E-11-1.02787872E+04 1.45722395E+01-1.30831522E+04    4
CH3CHCHCHO        T 5/92C   4H   6O   1    0G   298.150  3000.0    1000.0      1
 1.98794540E+01-2.09130550E-02 4.45360508E-05-2.60374870E-08 4.86836120E-12    2
-1.95278768E+04-6.87200320E+01-1.55577660E+00 4.09640630E-02-1.69868810E-05    3
-6.00928140E-18 2.31368530E-21-1.41394920E+04 3.74707580E+01-1.29340710E+04    4
C4H4O             T03/97C   4H   4O   1    0G   200.000  6000.0    1000.0      1
 9.38935003E+00 1.40291241E-02-5.07755110E-06 8.24137332E-10-4.95319963E-14    2
-8.68241814E+03-2.79162920E+01 8.47469463E-01 1.31773796E-02 5.99735901E-05    3
-9.71562904E-08 4.22733796E-11-5.36785445E+03 2.14945172E+01-4.17166616E+03    4
H2CC              L12/89H   2C   2    0    0G   200.000  6000.000  1000.000    1
 0.42780340E+01 0.47562804E-02-0.16301009E-05 0.25462806E-09-0.14886379E-13    2
 0.48316688E+05 0.64023701E+00 0.32815483E+01 0.69764791E-02-0.23855244E-05    3
-0.12104432E-08 0.98189545E-12 0.48621794E+05 0.59203910E+01 0.49887266E+05    4
H2C4O             120189H   2C   4O   1     G  0300.00   4000.00  1000.00      1
 0.01026888E+03 0.04896164E-01-0.04885081E-05-0.02708566E-08 0.05107013E-12    2
 0.02346903E+06-0.02815985E+03 0.04810971E+02 0.01313999E+00 0.09865073E-05    3
-0.06120720E-07 0.01640003E-10 0.02545803E+06 0.02113424E+02                   4
C6H2              P 1/93C   6H   2    0    0G   300.000  3000.00  1000.00      1
 0.13226281E+02 0.73904302E-02-0.22715381E-05 0.25875217E-09-0.55356741E-14    2
 0.80565258E+05-0.41201176E+02-0.15932624E+01 0.80530145E-01-0.14800649E-03    3
 0.13300031E-06-0.45332313E-10 0.83273227E+05 0.27980873E+02                   4
C6H3              H6W/94C   6H   3    0    0G   300.000  3000.00  1000.00      1
 0.58188343E+01 0.27933408E-01-0.17825427E-04 0.53702536E-08-0.61707627E-12    2
 0.85188250E+05-0.92147827E+00 0.11790619E+01 0.55547360E-01-0.73076168E-04    3
 0.52076736E-07-0.15046964E-10 0.85647312E+05 0.19179199E+02                   4
L-C6H4            H6W/94C   6H   4    0    0G   300.000  3000.00  1000.00      1
 0.12715182E+02 0.13839662E-01-0.43765440E-05 0.31541636E-09 0.46619026E-13    2
 0.57031148E+05-0.39464600E+02 0.29590225E+00 0.58053318E-01-0.67766756E-04    3
 0.43376762E-07-0.11418864E-10 0.60001371E+05 0.22318970E+02                   4
C-C6H4            H6W/94C   6H   4    0    0G   300.000  3000.00  1000.00      1
 0.13849209E+02 0.78807920E-02 0.18243836E-05-0.21169166E-08 0.37459977E-12    2
 0.47446340E+05-0.50404953E+02-0.30991268E+01 0.54030564E-01-0.40839004E-04    3
 0.10738837E-07 0.98078490E-12 0.52205711E+05 0.37415207E+02                   4
C6H5OH            L 4/84C   6H   6O   1    0G   300.000  5000.000 1000.        1
 0.14912073E+02 0.18378135E-01-0.61983128E-05 0.91983221E-09-0.49209565E-13    2
-0.18375199E+05-0.55924103E+02-0.16956539E+01 0.52271299E-01-0.72024050E-05    3
-0.35859603E-07 0.20449073E-10-0.13284121E+05 0.32542160E+02-0.11594207E+05    4
C6H5O             T05/02C   6H   5O   1    0G   200.000  6000.000 1000.        1
 1.37221720E+01 1.74688771E-02-6.35504520E-06 1.03492308E-09-6.23410504E-14    2
 2.87274751E+02-4.88181680E+01-4.66204455E-01 4.13443975E-02 1.32412991E-05    3
-5.72872769E-08 2.89763707E-11 4.77858391E+03 2.76990274E+01 6.49467016E+03    4
P-C6H4O2          AK0405C   6H   4O   2    0G   270.000  3000.000 1370.00      1
 1.23423732E+01 2.40612690E-02-1.16565184E-05 2.71393504E-09-2.47643065E-13    2
-2.06185312E+04-4.08244024E+01-2.43170113E+00 6.87937608E-02-6.41382837E-05    3
 3.08126855E-08-5.99832072E-12-1.65696994E+04 3.48309430E+01                   4
P-C6H3O2          AK0505C   6H   3O   2    0G   270.000  3000.000 1290.00      1
 1.22963699E+01 2.15055142E-02-1.07516136E-05 2.57528163E-09-2.41023652E-13    2
 1.15428998E+04-3.72584002E+01-1.57852347E+00 6.55376473E-02-6.50308721E-05    3
 3.32026554E-08-6.86665555E-12 1.51750093E+04 3.31518638E+01                   4
O-C6H4O2          AK0405C   6H   4O   2    0G   270.000  3000.000 1370.00      1
 1.23614349E+01 2.40491397E-02-1.16529057E-05 2.71332785E-09-2.47593219E-13    2
-1.67079717E+04-4.00310857E+01-2.36179712E+00 6.86058343E-02-6.39129516E-05    3
 3.06903009E-08-5.97357785E-12-1.26704431E+04 3.53724482E+01                   4
C5H5             TAK0505C   5H   5    0    0G   298.150  3500.000  969.35      1
 1.33675715E+00 3.24793912E-02-1.67587774E-05 4.03514137E-09-3.70739036E-13    2
 3.00730524E+04 1.60315806E+01-3.97555452E+00 7.41370991E-02-1.11803345E-04    3
 9.04628776E-08-2.80999747E-11 3.01769405E+04 3.67153636E+01                   4
C5H6              T 1/90C   5H   6    0    0G   200.000  6000.000 1000.        1
 0.99757848E+01 0.18905543E-01-0.68411461E-05 0.11099340E-08-0.66680236E-13    2
 0.11081693E+05-0.32209454E+02 0.86108957E+00 0.14804031E-01 0.72108895E-04    3
-0.11338055E-06 0.48689972E-10 0.14801755E+05 0.21353453E+02 0.16152485E+05    4
C5H5OH     5/ 2/91 THE.MC   5H   6O   1    0G   300.000  5000.000 1398.000     1
 1.53433477E+01 1.50754059E-02-5.13553582E-06 7.95807816E-10-4.61311517E-14    2
-1.19645453E+04-5.85204430E+01-4.26822012E+00 6.62446749E-02-5.68494038E-05    3
 2.46858526E-08-4.26820696E-12-5.75581338E+03 4.47962850E+01                   4
C5H4O             T 8/99C   5H   4O   1    0G   200.000  6000.000 1000.        1
 1.00806824E+01 1.61143465E-02-5.83314509E-06 9.46759320E-10-5.68972206E-14    2
 1.94364771E+03-2.94521623E+01 2.64576497E-01 3.34873827E-02 1.67738470E-06    3
-2.96207455E-08 1.54431476E-11 5.11159287E+03 2.35409513E+01 6.64245999E+03    4
C5H5O      5/16/90 THERMC   5H   5O   1    0G   300.000  5000.000 1392.000     1
 1.48322894E+01 1.40483376E-02-4.92302051E-06 7.77041219E-10-4.56103939E-14    2
 1.45523665E+04-5.73228191E+01-2.83112840E+00 5.67277287E-02-4.44757303E-05    3
 1.74924447E-08-2.76004847E-12 2.04992154E+04 3.69634411E+01                   4
C5H4OH            T 8/99C   5H   5O   1    0G   200.000  6000.000 1000.        1
 1.33741248E+01 1.51996469E-02-5.45685046E-06 8.80944866E-10-5.27493258E-14    2
 2.20358027E+03-4.59569069E+01-1.28398054E+00 4.90298511E-02-1.35844414E-05    3
-2.92983743E-08 1.90820619E-11 6.37364803E+03 3.08073591E+01 8.00114499E+03    4
C6H5OO     3/26/ 9 THERMC   6H   5O   2    0G   300.000  5000.000 1403.000     1
 1.67078262E+01 1.62326229E-02-5.47969630E-06 8.43510060E-10-4.86562431E-14    2
 8.14242915E+03-6.08346973E+01-2.99164672E+00 7.03857150E-02-6.34400574E-05    3
 2.91548920E-08-5.30706938E-12 1.41320240E+04 4.20142955E+01                   4
C6H5OOH    3/26/ 9 THERMC   6H   6O   2    0G   300.000  5000.000 1404.000     1
 1.92317474E+01 1.63154699E-02-5.53448904E-06 8.55059974E-10-4.94583790E-14    2
-1.01971012E+04-7.61674471E+01-4.03105975E+00 7.96101888E-02-7.21655013E-05    3
 3.27610696E-08-5.85584239E-12-3.10973017E+03 4.54324978E+01                   4
C6H4OH     4/ 9/ 9 THERMC   6H   5O   1    0G   300.000  5000.000 1402.000     1
 1.73187560E+01 1.36366984E-02-4.68316332E-06 7.29071204E-10-4.23805358E-14    2
 1.14990276E+04-6.89986593E+01-5.99875435E+00 8.59063379E-02-9.12525636E-05    3
 4.72275890E-08-9.35576749E-12 1.78621926E+04 4.99931427E+01                   4
HOC6H4OH   4/ 9/ 9 THERMC   6H   6O   2    0G   300.000  5000.000 1405.000     1
 2.31394847E+01 1.31873680E-02-4.49072464E-06 6.95268891E-10-4.02643108E-14    2
-4.25885990E+04-1.02692352E+02-8.68529064E+00 1.17282933E-01-1.33754802E-04    3
 7.16697462E-08-1.44385730E-11-3.44903827E+04 5.77087257E+01                   4
OC6H4OH    4/ 9/ 9 THERMC   6H   5O   2    0G   300.000  5000.000 1403.000     1
 2.22718210E+01 1.21038561E-02-4.18429526E-06 6.54475399E-10-3.81746504E-14    2
-2.34827539E+04-9.61035467E+01-8.02205657E+00 1.09403210E-01-1.23489276E-04    3
 6.56286805E-08-1.31527870E-11-1.55949156E+04 5.72175202E+01                   4
P-OC6H5OJ  WKM          C   6O   2H   5    0G   300.000  5000.000 1400.000     1
 1.82799770E+01 1.59280974E-02-5.50765220E-06 8.61649836E-10-5.02677539E-14    2
-6.25907994E+01-7.25809444E+01-3.29683290E+00 7.27365977E-02-6.36158220E-05    3
 2.80683553E-08-4.92279426E-12 6.73402222E+03 4.09349895E+01                   4
O-OC6H5OJ  WKM          C   6O   2H   5    0G   300.000  5000.000 1400.000     1
 1.84625733E+01 1.57607263E-02-5.44671499E-06 8.51765760E-10-4.96759541E-14    2
-1.72770226E+02-7.28742484E+01-2.65459198E+00 7.17179095E-02-6.31552372E-05    3
 2.81132946E-08-4.97463333E-12 6.45283150E+03 3.81123139E+01                   4
C#CC*CCJ           GLAR C   5H   5    0    0G   300.000  5000.000 1396.000     1
 1.41230912E+01 1.14233190E-02-3.95851276E-06 6.20128961E-10-3.62097887E-14    2
 4.25158384E+04-5.02942871E+01-6.16143558E-01 5.06466579E-02-4.48561743E-05    3
 2.02459419E-08-3.64542145E-12 4.71532377E+04 2.71623299E+01                   4
C5H6-L     2/ 5/ 9 THERMC   5H   6    0    0G   300.000  5000.000 1372.000     1
 1.29600892E+01 1.48953758E-02-5.23622902E-06 8.27916389E-10-4.86464523E-14    2
 2.38180800E+04-4.25312093E+01 3.58448213E+00 3.24459626E-02-1.70150991E-05    3
 4.22715914E-09-4.18452556E-13 2.76514681E+04 9.60644208E+00                   4
CJ*CC*CC*O 2/ 5/ 9 THERMC   5H   5O   1    0G   300.000  5000.000 1396.000     1
 1.62360823E+01 1.18297101E-02-4.11454219E-06 6.46026823E-10-3.77767639E-14    2
 1.93499885E+04-5.83498817E+01-5.06628841E-01 6.04671965E-02-5.97396749E-05    3
 2.96804228E-08-5.76240010E-12 2.42765544E+04 2.82994148E+01                   4
C*CC*CCJ*O 2/ 5/ 9 THERMC   5H   5O   1    0G   300.000  5000.000 1399.000     1
 1.53178248E+01 1.27352911E-02-4.35882964E-06 6.76912763E-10-3.92771371E-14    2
 7.60582726E+03-5.43599625E+01-2.18492198E-01 5.92100223E-02-5.89241174E-05    3
 2.97411920E-08-5.85244770E-12 1.20600764E+04 2.55968530E+01                   4
CJ*CC*O    4/ 8/94 THERMC   3H   3O   1    0G   300.000  5000.000 1402.000     1
 1.07482537E+01 6.19822688E-03-2.06130981E-06 3.14418872E-10-1.80309517E-14    2
 1.51410162E+04-3.01266033E+01 1.46654466E+00 3.23390476E-02-3.05588208E-05    3
 1.44081861E-08-2.65600505E-12 1.78850058E+04 1.80850321E+01                   4
C5H3O            TAK0905C   5H   3O   1    0G   300.000  3500.000 1500.00      1
 1.19961781E+01 1.34287065E-02-5.90045309E-06 1.22553862E-09-9.86114716E-14    2
 2.89592010E+04-4.07548249E+01-3.03242604E+00 5.43937201E-02-4.95018348E-05    3
 2.25523751E-08-4.10727920E-12 3.35644081E+04 3.78374823E+01                   4
C5H7       1/22/ 9 WKM  C   5H   7    0    0G   300.000  5000.000 1377.000     1
 1.36630213E+01 1.68061358E-02-5.98746539E-06 9.55341072E-10-5.64951981E-14    2
 1.27238941E+04-5.46331286E+01-6.75118368E+00 6.06461693E-02-4.01260152E-05    3
 1.22051562E-08-1.33459844E-12 2.01365277E+04 5.62694938E+01                   4
OC5H7O     1/22/ 9 WKM  C   5H   7O   2    0G   300.000  5000.000 1375.000     1
 1.65416953E+01 1.86677673E-02-6.44836048E-06 1.00787611E-09-5.87521858E-14    2
-2.82017168E+04-5.47258181E+01 4.88394767E+00 4.03401300E-02-1.97774150E-05    3
 3.68903501E-09-3.40202384E-14-2.35295942E+04 9.97070337E+00                   4
C*CCJC*COH 10/6/95 Z&B  C   5H   7O   1    0G   300.000  5000.000 1397.000     1
 1.67465815E+01 1.58357240E-02-5.44954706E-06 8.49881387E-10-4.94743246E-14    2
-4.30972870E+03-6.19378748E+01-2.91175436E+00 6.69362484E-02-5.71603047E-05    3
 2.48753749E-08-4.33243894E-12 1.96441523E+03 4.17454344E+01                   4
C*CC*CCJ           Z&B  C   5H   7    0    0G   300.000  5000.000 1386.000     1
 1.47302883E+01 1.59030900E-02-5.57729508E-06 8.80604825E-10-5.16963733E-14    2
 1.74050791E+04-5.42670706E+01-1.60087476E+00 5.38764703E-02-3.96302225E-05    3
 1.49599474E-08-2.31995284E-12 2.31199746E+04 3.35492960E+01                   4
C*CC*CC    3/1/95  Z&B  C   5H   8    0    0G   300.000  5000.000 1395.000     1
 1.41303131E+01 1.81877961E-02-6.19208788E-06 9.58333792E-10-5.54785472E-14    2
 2.25907168E+03-5.11705577E+01-1.19376866E+00 5.65474329E-02-4.39472481E-05    3
 1.82341266E-08-3.12226566E-12 7.36084709E+03 3.02808980E+01                   4
C*CC*CCOH  1/23/ 9 WKM  C   5H   8O   1    0G   300.000  5000.000 1396.000     1
 1.63079670E+01 1.79957763E-02-6.03115896E-06 9.23992259E-10-5.31254053E-14    2
-1.58204603E+04-5.84137244E+01-5.31488384E-01 6.06983915E-02-4.81499862E-05    3
 2.00308244E-08-3.38987282E-12-1.03301302E+04 3.07961436E+01                   4
C*CCJC*O           Z&B  C   4H   5O   1    0G   300.000  5000.000 1385.000     1
 1.22833215E+01 1.26428506E-02-4.31034879E-06 6.68415867E-10-3.87693974E-14    2
 1.86818728E+03-3.84807909E+01-4.83886977E-01 4.23431670E-02-3.05389089E-05    3
 1.11441978E-08-1.63863920E-12 6.28635090E+03 3.00860103E+01                   4
OC4H6O     1/23/ 9 WKM  C   4H   6O   2    0G   300.000  5000.000 1382.000     1
 1.41894774E+01 1.53345510E-02-5.24594862E-06 8.14655154E-10-4.72759368E-14    2
-4.10001835E+04-4.43771751E+01 4.21628848E+00 3.57422725E-02-2.04226185E-05    3
 5.63821367E-09-5.88888993E-13-3.72055911E+04 1.02814620E+01                   4
OC4H5O     1/23/ 9 WKM  C   4H   5O   2    0G   300.000  5000.000 1388.000     1
 1.32138775E+01 1.37339051E-02-4.62639517E-06 7.10941370E-10-4.09538499E-14    2
-2.16535271E+04-3.64185255E+01 4.60550978E+00 3.30498712E-02-2.13102363E-05    3
 7.37021089E-09-1.08289438E-12-1.85460831E+04 1.01599453E+01                   4
HOC*CC*O   1/26/ 9 WKM  C   3H   4O   2    0G   300.000  5000.000 1413.000     1
 1.66505478E+01 6.11745137E-03-2.09080785E-06 3.24985683E-10-1.88875073E-14    2
-3.82179939E+04-6.36794754E+01-2.01837189E+00 6.26539783E-02-6.73359280E-05    3
 3.39430425E-08-6.48917648E-12-3.31367523E+04 3.18162860E+01                   4
HOC*CCJ*O  1/26/ 9 WKM  C   3H   3O   2    0G   300.000  5000.000 1414.000     1
 1.52720985E+01 5.02586331E-03-1.68408578E-06 2.58390706E-10-1.48849424E-14    2
-1.98506828E+04-5.54641734E+01 6.07270082E-01 4.96011303E-02-5.32300885E-05    3
 2.68392951E-08-5.13094510E-12-1.58814562E+04 1.94817133E+01                   4
C2H2OH                  H   3C   2O   1    0G    300.00   5000.00 1000.00      1
 6.81339897E+00 8.05827723E-03-3.11728612E-06 5.54590896E-10-3.71804255E-14    2
 1.31583034E+04-1.09863525E+01 5.62397968E-01 2.64598620E-02-2.28453705E-05    3
 9.14478695E-09-1.06711936E-12 1.48374643E+04 2.10439544E+01                   4
O2CCHOOJ           Z&B  C   2H   1O   4    0G   300.000  5000.000 1682.000     1
 1.09910849E+01 7.46985861E-03-2.75568271E-06 4.51353051E-10-2.72108652E-14    2
-3.51335323E+04-2.11652231E+01 8.91497688E+00 8.60571847E-03 5.24416766E-07    3
-2.79301331E-09 7.62963051E-13-3.40867754E+04-8.72978273E+00                   4
HCOH              MAR94 C   1H   2O   1    0G   300.     5000.    1398.        1
 9.18749272E+00 1.52011152E-03-6.27603516E-07 1.09727989E-10-6.89655128E-15    2
 7.81364593E+03-2.73434214E+01-2.82157421E+00 3.57331702E-02-3.80861580E-05    3
 1.86205951E-08-3.45957838E-12 1.12956672E+04 3.48487757E+01                   4
C2H3OH     2/ 3/ 9 THERMC   2H   4O   1    0G   300.000  5000.000 1410.000     1
 8.32598158E+00 8.03387281E-03-2.63928405E-06 3.98410726E-10-2.26551155E-14    2
-1.83221436E+04-2.02080305E+01-1.27972260E-01 3.38506073E-02-3.30644935E-05    3
 1.64858739E-08-3.19935455E-12-1.59914544E+04 2.30438601E+01                   4
O2CH2CHO          BOZ_03C   2H   3O   3    0G   300.000  5000.000 1393.000     1
 1.11807543E+01 9.14479256E-03-3.15089833E-06 4.91944238E-10-2.86639180E-14    2
-1.55790331E+04-2.87892740E+01-1.29465843E+00 4.44936393E-02-4.26577074E-05    3
 2.07391950E-08-3.96828771E-12-1.18275628E+04 3.60778797E+01                   4
HO2CH2CO          BOZ_03C   2H   3O   3    0G   300.000  5000.000 1386.000     1
 1.04146322E+01 1.12680116E-02-5.17494839E-06 1.00333285E-09-6.68165911E-14    2
-1.40955672E+04-2.27894400E+01 2.22681686E+00 3.56781380E-02-3.26401909E-05    3
 1.47651988E-08-2.64794380E-12-1.18735095E+04 1.91581197E+01                   4
END


