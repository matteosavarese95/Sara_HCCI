THERMO ALL
300.  1000.  5000.
AR                G 5/97AR  1  0    0      0G   200.000  6000.00  1000.00      1
+2.50000000E+00+0.00000000E+00+0.00000000E+00+0.00000000E+00+0.00000000E+00    2
-7.45375000E+02+4.37967491E+00+2.50000000E+00+0.00000000E+00+0.00000000E+00    3
+0.00000000E+00+0.00000000E+00-7.45375000E+02+4.37967491E+00+0.00000000E+00    4
N2                G 8/02N   2    0    0    0G   200.000  6000.00  1000.00      1
+2.95257637E+00+1.39690040E-03-4.92631603E-07+7.86010195E-11-4.60755204E-15    2
-9.23948688E+02+5.87188762E+00+3.53100528E+00-1.23660988E-04-5.02999433E-07    3
+2.43530612E-09-1.40881235E-12-1.04697628E+03+2.96747038E+00+0.00000000E+00    4
HE                G 5/97HE 1    0    0    0 G   200.000  6000.00  1000.00      1
+2.50000000E+00+0.00000000E+00+0.00000000E+00+0.00000000E+00+0.00000000E+00    2
-7.45375000E+02+9.28723974E-01+2.50000000E+00+0.00000000E+00+0.00000000E+00    3
+0.00000000E+00+0.00000000E+00-7.45375000E+02+9.28723974E-01+0.00000000E+00    4
H2                TPIS78H   2    0    0    0G   200.000  6000.00  1000.00      1
+2.93286575E+00+8.26608026E-04-1.46402364E-07+1.54100414E-11-6.88804800E-16    2
-8.13065581E+02-1.02432865E+00+2.34433112E+00+7.98052075E-03-1.94781510E-05    3
+2.01572094E-08-7.37611761E-12-9.17935173E+02+6.83010238E-01+0.00000000E+00    4
H                 L 6/94H   1    0    0    0G   200.000  6000.00  1000.00      1
+2.50000000E+00+0.00000000E+00+0.00000000E+00+0.00000000E+00+0.00000000E+00    2
+2.54736600E+04-4.46682850E-01+2.50000000E+00+0.00000000E+00+0.00000000E+00    3
+0.00000000E+00+0.00000000E+00+2.54736600E+04-4.46682850E-01+2.62190350E+04    4
O2                RUS 89O   2    0    0    0G   200.000  6000.00  1000.00      1
+3.66096065E+00+6.56365811E-04-1.41149627E-07+2.05797935E-11-1.29913436E-15    2
-1.21597718E+03+3.41536279E+00+3.78245636E+00-2.99673416E-03+9.84730201E-06    3
-9.68129509E-09+3.24372837E-12-1.06394356E+03+3.65767573E+00+0.00000000E+00    4
O                 L 1/90O   1    0    0    0G   200.000  6000.00  1000.00      1
+2.54363697E+00-2.73162486E-05-4.19029520E-09+4.95481845E-12-4.79553694E-16    2
+2.92260120E+04+4.92229457E+00+3.16826710E+00-3.27931884E-03+6.64306396E-06    3
-6.12806624E-09+2.11265971E-12+2.91222592E+04+2.05193346E+00+2.99687009E+04    4
H2O               L 5/89H   2 O  1    0    0G   200.000  6000.00  1000.00      1
+2.67703890E+00+2.97318160E-03-7.73768890E-07+9.44335140E-11-4.26899910E-15    2
-2.98858940E+04+6.88255000E+00+4.19863520E+00-2.03640170E-03+6.52034160E-06    3
-5.48792690E-09+1.77196800E-12-3.02937260E+04-8.49009010E-01-2.90848170E+04    4
OH                IU3/03O   1 H  1    0    0G   200.000  6000.00  1000.00      1
+2.83853033E+00+1.10741289E-03-2.94000209E-07+4.20698729E-11-2.42289890E-15    2
+3.69780808E+03+5.84494652E+00+3.99198424E+00-2.40106655E-03+4.61664033E-06    3
-3.87916306E-09+1.36319502E-12+3.36889836E+03-1.03998477E-01+4.48613328E+03    4
OHV       11/13/18 THERMC   0H   1O   1    0G   300.000  5000.000 1710.000     1
 2.85376040E+00 1.02994334E-03-2.32666477E-07 1.93750704E-11-3.15759847E-16    2
 5.03225473E+04 5.76240468E+00 3.41896226E+00 3.19255801E-04-3.08292717E-07    3
 3.64407494E-10-1.00195479E-13 5.00756946E+04 2.51917016E+00                   4
H2O2              T 8/03H   2O   2    0    0G   200.000  6000.00  1000.00      1
+4.57977305E+00+4.05326003E-03-1.29844730E-06+1.98211400E-10-1.13968792E-14    2
-1.80071775E+04+6.64970694E-01+4.31515149E+00-8.47390622E-04+1.76404323E-05    3
-2.26762944E-08+9.08950158E-12-1.77067437E+04+3.27373319E+00-1.63425145E+04    4
HO2               T 1/09H   1O   2    0    0G   200.000  5000.00  1000.00      1
+4.17228741E+00+1.88117627E-03-3.46277286E-07+1.94657549E-11+1.76256905E-16    2
+3.10206839E+01+2.95767672E+00+4.30179807E+00-4.74912097E-03+2.11582905E-05    3
-2.42763914E-08+9.29225225E-12+2.64018485E+02+3.71666220E+00+1.47886045E+03    4
CO                RUS 79C   1O   1    0    0G   200.000  6000.00  1000.00      1
+3.04848590E+00+1.35172810E-03-4.85794050E-07+7.88536440E-11-4.69807460E-15    2
-1.42661170E+04+6.01709770E+00+3.57953350E+00-6.10353690E-04+1.01681430E-06    3
+9.07005860E-10-9.04424490E-13-1.43440860E+04+3.50840930E+00-1.32936280E+04    4
CO2               L 7/88C   1O   2    0    0G   200.000  6000.00  1000.00      1
+4.63651110E+00+2.74145690E-03-9.95897590E-07+1.60386660E-10-9.16198570E-15    2
-4.90249040E+04-1.93489550E+00+2.35681300E+00+8.98412990E-03-7.12206320E-06    3
+2.45730080E-09-1.42885480E-13-4.83719710E+04+9.90090350E+00-4.73281050E+04    4
HOCO              T05/06H  1 C  1 O  2    0 G   200.000  6000.00   1000.00     1
+5.39206152E+00+4.11221455E-03-1.48194900E-06+2.39875460E-10-1.43903104E-14    2
-2.38606717E+04-2.23529091E+00+2.92207919E+00+7.62453859E-03+3.29884437E-06    3
-1.07135205E-08+5.11587057E-12-2.30281524E+04+1.12925886E+01-2.18076591E+04    4
CH4               G 8/99C  1 H  4    0    0 G   200.000  6000.00  1000.00      1
+1.65326226E+00+1.00263099E-02-3.31661238E-06+5.36483138E-10-3.14696758E-14    2
-1.00095936E+04+9.90506283E+00+5.14911468E+00-1.36622009E-02+4.91453921E-05    3
-4.84246767E-08+1.66603441E-11-1.02465983E+04-4.63848842E+00-8.97226656E+03    4
CH3               IU0702C  1 H  3    0    0 G   200.000  6000.00  1000.00      1
+2.97812060E+00+5.79785200E-03-1.97558000E-06+3.07297900E-10-1.79174160E-14    2
+1.65095130E+04+4.72247990E+00+3.65717970E+00+2.12659790E-03+5.45838830E-06    3
-6.61810030E-09+2.46570740E-12+1.64227160E+04+1.67353540E+00+1.76439350E+04    4
CH2               IU3/03C  1 H  2    0    0 G   200.000  6000.00  1000.00      1
+3.14631886E+00+3.03671259E-03-9.96474439E-07+1.50483580E-10-8.57335515E-15    2
+4.60412605E+04+4.72341711E+00+3.71757846E+00+1.27391260E-03+2.17347251E-06    3
-3.48858500E-09+1.65208866E-12+4.58723866E+04+1.75297945E+00+4.70504920E+04    4
CH2(S)            IU6/03C  1 H  2    0    0 G   200.000  6000.00  1000.00      1
+3.13501686E+00+2.89593926E-03-8.16668090E-07+1.13572697E-10-6.36262835E-15    2
+5.05040504E+04+4.06030621E+00+4.19331325E+00-2.33105184E-03+8.15676451E-06    3
-6.62985981E-09+1.93233199E-12+5.03662246E+04-7.46734310E-01+5.15727280E+04    4
C                 L 7/88C   1     0    0   0G   200.000  6000.00  1000.00      1
+2.60558300E+00-1.95934340E-04+1.06737220E-07-1.64239400E-11+8.18705800E-16    2
+8.54117420E+04+4.19238680E+00+2.55423950E+00-3.21537720E-04+7.33792230E-07    3
-7.32234870E-10+2.66521440E-13+8.54426810E+04+4.53130850E+00+8.61950970E+04    4
CH                IU3/03C  1 H  1    0    0 G   200.000  6000.00  1000.00      1
+2.52093690E+00+1.76536390E-03-4.61476600E-07+5.92896750E-11-3.34745010E-15    2
+7.09467690E+04+7.40518290E+00+3.48975830E+00+3.24321600E-04-1.68997510E-06    3
+3.16284200E-09-1.40618030E-12+7.06126460E+04+2.08428410E+00+7.16581880E+04    4
CHV       11/13/18 THERMC   1H   1O   0    0G   300.000  5000.000 1365.000     1
 2.21703785E+00 2.15314038E-03-5.71569209E-07 6.54441183E-11-2.66374894E-15    2
 1.04414085E+05 9.18247549E+00 3.50775836E+00-4.57470019E-04 1.32602633E-06    3
-5.14213760E-10 5.82219975E-14 1.03920991E+05 2.09911232E+00                   4
CH3O2H            A 7/05C  1 H  4 O  2    0 G   200.000  6000.00  1000.00      1
+7.76538058E+00+8.61499712E-03-2.98006935E-06+4.68638071E-10-2.75339255E-14    2
-1.82979984E+04-1.43992663E+01+2.90540897E+00+1.74994735E-02+5.28243630E-06    3
-2.52827275E-08+1.34368212E-11-1.68894632E+04+1.13741987E+01-1.52423685E+04    4
CH3O2                   H   3C   1O   2    0G   300.000  5000.000 1374.000     1
+6.47970487E+00+7.44401080E-03-2.52348555E-06+3.89577296E-10-2.25182399E-14    2
-1.56285441E+03-8.19477074E+00+1.97339205E+00+1.53542340E-02-6.37314891E-06    3
+3.19930565E-10+2.82193915E-13+2.54278835E+02+1.69194215E+01+0.00000000E+00    4
CH2O2H     9/ 1/12      C   1H   3O   2    0G   300.000  5000.000 1410.000     2
+9.24697852E+00+4.60845541E-03-1.53501472E-06+2.34434830E-10-1.34573106E-14    2
+4.11529953E+03-2.11503248E+01+2.88976454E+00+2.09465776E-02-1.75190772E-05    3
+7.27819787E-09-1.18912344E-12+6.12390620E+03+1.23802076E+01+0.00000000E+00    4
CH3OH             T06/02C   1H  4 O  1    0 G   200.000  6000.00  1000.00      1
+3.52726795E+00+1.03178783E-02-3.62892944E-06+5.77448016E-10-3.42182632E-14    2
-2.60028834E+04+5.16758693E+00+5.65851051E+00-1.62983419E-02+6.91938156E-05    3
-7.58372926E-08+2.80427550E-11-2.56119736E+04-8.97330508E-01-2.41746056E+04    4
CH3O              IU1/03C  1 H  3 O  1    0 G   200.000  6000.00  1000.00      1
+4.75779238E+00+7.44142474E-03-2.69705176E-06+4.38090504E-10-2.63537098E-14    2
+3.78111940E+02-1.96680028E+00+3.71180502E+00-2.80463306E-03+3.76550971E-05    3
-4.73072089E-08+1.86588420E-11+1.29569760E+03+6.57240864E+00+2.52571660E+03    4
CH2OH             IU2/03C  1 H  3 O  1    0 G   200.000  6000.00   1000.00     1
+5.09314370E+00+5.94761260E-03-2.06497460E-06+3.23008173E-10-1.88125902E-14    2
-4.03409640E+03-1.84691493E+00+4.47834367E+00-1.35070310E-03+2.78484980E-05    3
-3.64869060E-08+1.47907450E-11-3.50072890E+03+3.30913500E+00-2.04462770E+03    4
CH2O              T 5/11H   2C   1O   1    0G   200.000  6000.00  1000.00      1
+3.16952665E+00+6.19320560E-03-2.25056366E-06+3.65975660E-10-2.20149458E-14    2
-1.45486831E+04+6.04207898E+00+4.79372312E+00-9.90833322E-03+3.73219990E-05    3
-3.79285237E-08+1.31772641E-11-1.43791953E+04+6.02798058E-01-1.31293365E+04    4
HCO               T 5/03C  1 H  1 O  1    0 G   200.000  6000.00  1000.00      1
+3.92001542E+00+2.52279324E-03-6.71004164E-07+1.05615948E-10-7.43798261E-15    2
+3.65342928E+03+3.58077056E+00+4.23754610E+00-3.32075257E-03+1.40030264E-05    3
-1.34239995E-08+4.37416208E-12+3.87241185E+03+3.30834869E+00+5.08749163E+03    4
HCOH              MAR94 C   1H   2O   1    0G   300.     5000.    1398.        1
+9.18749272E+00+1.52011152E-03-6.27603516E-07+1.09727989E-10-6.89655128E-15    2
+7.81364593E+03-2.73434214E+01-2.82157421E+00+3.57331702E-02-3.80861580E-05    3
+1.86205951E-08-3.45957838E-12+1.12956672E+04+3.48487757E+01+0.00000000E+00    4
HO2CHO     6/26/95 THERMC   1H   2O   3    0G   300.000  5000.000 1378.00      2
+9.87503878E+00+4.64663708E-03-1.67230522E-06+2.68624413E-10-1.59595232E-14    2
-3.80502496E+04-2.24939155E+01+2.42464726E+00+2.19706380E-02-1.68705546E-05    3
+6.25612194E-09-9.11645843E-13-3.54828006E+04+1.75027796E+01+0.00000000E+00    4
HOCH2O2H   9/ 1/12      C   1H   4O   3    0G   300.000  5000.000 1398.000     2
+1.24531886E+01+7.18221110E-03-2.47029548E-06+3.85611737E-10-2.24774193E-14    2
-4.24862928E+04-3.58745197E+01+5.35189713E-01+3.73266553E-02-3.15299511E-05    3
+1.30352583E-08-2.11473264E-12-3.86609415E+04+2.71776082E+01+0.00000000E+00    4
HOCH2O2    9/ 1/12      C   1H   3O   3    0G   300.000  5000.000 1377.000     2
+1.16406115E+01+5.72826040E-03-2.05362036E-06+3.29070695E-10-1.95188360E-14    2
-2.53505769E+04-3.07332064E+01+2.82068616E+00+2.47857094E-02-1.66186399E-05    3
+4.79633095E-09-4.28087766E-13-2.22077036E+04+1.70599803E+01+0.00000000E+00    4
OCH2O2H    7/21/14 THERMC   1H   3O   3    0G   300.000  5000.000 1418.000     3
+1.29622491E+01+4.21948855E-03-1.54275194E-06+2.50413077E-10-1.49855537E-14    2
-1.81326406E+04-3.87016356E+01+4.46349361E-01+3.63049606E-02-3.26130978E-05    3
+1.37050551E-08-2.20872791E-12-1.41972598E+04+2.72960376E+01+0.00000000E+00    4
HOCH2O     2/16/99 THERMC   1H   3O   2    0G   300.000  5000.000 1452.000     1
+6.39521515E+00+7.43673043E-03-2.50422354E-06+3.84879712E-10-2.21778689E-14    2
-2.41108840E+04-6.63865583E+00+4.11183145E+00+7.53850697E-03+3.77337370E-06    3
-5.38746005E-09+1.45615887E-12-2.28023001E+04+7.46807254E+00+0.00000000E+00    4
O2CHO      6/26/95 THERMC   1H   1O   3    0G   300.000  5000.000 1368.00      1
+7.24075139E+00+4.63312951E-03-1.63693995E-06+2.59706693E-10-1.52964699E-14    2
-1.87027618E+04-6.49547212E+00+3.96059309E+00+1.06002279E-02-5.25713351E-06    3
+1.01716726E-09-2.87487602E-14-1.73599383E+04+1.17807483E+01+0.00000000E+00    4
HOCHO             L 8/88H   2C   1O   2    0G   200.000  6000.00  1000.00      1
+4.61383160E+00+6.44963640E-03-2.29082510E-06+3.67160470E-10-2.18736750E-14    2
-4.75148500E+04+8.47883830E-01+3.89836160E+00-3.55877950E-03+3.55205380E-05    3
-4.38499590E-08+1.71077690E-11-4.67706090E+04+7.34953970E+00-4.55312460E+04    4
OCHO              ATCT/AC  1 O  2 H  1    0 G   200.000  6000.000 1000.00      1
+4.14394211E+00+5.59738818E-03-1.99794019E-06+3.16179193E-10-1.85614483E-14    2
-1.72459887E+04+5.07778617E+00+4.68825921E+00-4.14871834E-03+2.55066010E-05    3
-2.84473900E-08+1.04422559E-11-1.69867041E+04+4.28426480E+00-1.55992356E+04    4
C2H6              G 8/88C   2H 6    0      0G   200.000  6000.00  1000.00      1
+4.04666411E+00+1.53538802E-02-5.47039485E-06+8.77826544E-10-5.23167531E-14    2
-1.24473499E+04-9.68698313E-01+4.29142572E+00-5.50154901E-03+5.99438458E-05    3
-7.08466469E-08+2.68685836E-11-1.15222056E+04+2.66678994E+00-1.00849652E+04    4
C2H5       8/ 4/ 4 THERMC   2H   5    0    0G   300.000  5000.000 1387.000     1
+5.88784390E+00+1.03076793E-02-3.46844396E-06+5.32499257E-10-3.06512651E-14    2
+1.15065499E+04-8.49651771E+00+1.32730217E+00+1.76656753E-02-6.14926558E-06    3
-3.01143466E-10+4.38617775E-13+1.34284028E+04+1.71789216E+01+0.00000000E+00    4
C2H5O2H    9/ 1/12      C   2H   6O   2    0G   300.000  5000.000 1390.000     3
+1.04823538E+01+1.34779879E-02-4.62179078E-06+7.18618519E-10-4.17307436E-14    2
-2.46578171E+04-2.84294243E+01+1.83755328E+00+3.38053586E-02-2.37548140E-05    3
+9.31974865E-09-1.58003428E-12-2.15814086E+04+1.80977584E+01+0.00000000E+00    4
C2H5O2     9/ 1/12      C   2H   5O   2    0G   300.000  5000.000 1389.000     2
+9.50282570E+00+1.20429839E-02-4.09491581E-06+6.33049241E-10-3.66133788E-14    2
-7.37069391E+03-2.21717130E+01+3.90351912E+00+2.22599212E-02-1.01610079E-05    3
+1.71709751E-09+1.88166738E-14-5.09654081E+03+8.98722750E+00+0.00000000E+00    4
C2H4       8/12/15      C   2H   4    0    0G   300.000  5000.000 1392.000     1
+5.07061289E+00+9.11140768E-03-3.10506692E-06+4.80733851E-10-2.78321396E-14    2
+3.66391217E+03-6.64501414E+00+4.81118223E-01+1.83778060E-02-9.99633565E-06    3
+2.73211039E-09-3.01837289E-13+5.44386648E+03+1.85867157E+01+0.00000000E+00    4
C2H3       8/12/15      C   2H   3    0    0G   300.000  5000.000 1400.000     1
+4.99675415E+00+6.55838271E-03-2.20921909E-06+3.39300272E-10-1.95316926E-14    2
+3.34604382E+04-3.01451097E+00+1.25545094E+00+1.57481597E-02-1.12218328E-05    3
+4.50915682E-09-7.74861577E-13+3.47435574E+04+1.69664043E+01+0.00000000E+00    4
CHOCHO                  C   2H   2O   2    0G   300.000  5000.000 1386.000     1
+9.75438561E+00+4.97645947E-03-1.74410483E-06+2.75586994E-10-1.61969892E-14    2
-2.95832896E+04-2.61878329E+01+1.88105120E+00+2.36386368E-02-1.83443295E-05    3
+6.84842963E-09-9.92733674E-13-2.69280190E+04+1.59154793E+01+0.00000000E+00    4
C2H3OOH    4/18/ 8 THERMC   2H   4O   2    0G   300.000  5000.000 1397.000     2
+1.15749951E+01+8.09909174E-03-2.81808668E-06+4.42697954E-10-2.58998042E-14    2
-8.84852664E+03-3.43859117E+01+1.35644398E+00+3.37002447E-02-2.75988500E-05    3
+1.14222854E-08-1.89488886E-12-5.49996692E+03+1.98354466E+01+0.00000000E+00    4
C2H3OO                  H   3C   2O   2     G   298.150  2000.000 1000.00      1
+6.04483828E+00+1.45511127E-02-7.50974622E-06+1.83488280E-09-1.66689681E-13    2
+1.01699244E+04-3.71144913E+00+1.09784776E+00+2.95333237E-02-2.27744360E-05    3
+7.20559155E-09-3.07929092E-13+1.13996101E+04+2.13563583E+01+0.00000000E+00    4
CHCHO                   H   2C   2O   1     G   298.150  2000.000 1000.00      1
+4.92632910E+00+9.71712147E-03-5.54855980E-06+1.53068537E-09-1.64742462E-13    2
+2.89499494E+04+5.27874677E-01+2.33256751E+00+1.62952986E-02-9.72052177E-06    3
+5.15124155E-10+1.03836514E-12+2.96585452E+04+1.39904923E+01+0.00000000E+00    4
C2H2              G 1/91C  2 H  2    0    0 G   200.000  6000.00  1000.00      1
+4.65878489E+00+4.88396667E-03-1.60828888E-06+2.46974544E-10-1.38605959E-14    2
+2.57594042E+04-3.99838194E+00+8.08679682E-01+2.33615762E-02-3.55172234E-05    3
+2.80152958E-08-8.50075165E-12+2.64289808E+04+1.39396761E+01+2.74459950E+04    4
C2H               T 5/10C  2 H  1    0    0 G   200.000  6000.00  1000.00      1
+3.66270248E+00+3.82492252E-03-1.36632500E-06+2.13455040E-10-1.23216848E-14    2
+6.71683790E+04+3.92205792E+00+2.89867676E+00+1.32988489E-02-2.80733327E-05    3
+2.89484755E-08-1.07502351E-11+6.70616050E+04+6.18547632E+00+6.83210436E+04    4
H2CC              L12/89H   2C   2    0    0G   200.000  6000.000  1000.000    1
+4.27803400E+00+4.75628040E-03-1.63010090E-06+2.54628060E-10-1.48863790E-14    2
+4.83166880E+04+6.40237010E-01+3.28154830E+00+6.97647910E-03-2.38552440E-06    3
-1.21044320E-09+9.81895450E-13+4.86217940E+04+5.92039100E+00+4.98872660E+04    4
C2H5OH     8/12/15      C   2H   6O   1    0G   300.000  5000.000 1402.000     2
+8.14483865E+00+1.28314052E-02-4.29052743E-06+6.55971721E-10-3.76506611E-14    2
-3.24005526E+04-1.86241126E+01+2.15805861E-01+2.95228396E-02-1.68271048E-05    3
+4.49484797E-09-4.02451543E-13-2.94851823E+04+2.45725052E+01+0.00000000E+00    4
C2H5O      8/12/15      C   2H   5O   1    0G   300.000  5000.000 1467.000     1
+8.19120635E+00+1.10391986E-02-3.75270536E-06+5.80275784E-10-3.35735146E-14    2
-5.66847208E+03-1.90131344E+01+2.90353584E+00+1.77256708E-02-2.69624757E-06    3
-3.45830533E-09+1.25224784E-12-3.28930290E+03+1.13545591E+01+0.00000000E+00    4
PC2H4OH    8/12/15      C   2H   5O   1    0G   300.000  5000.000 1395.000     2
+8.06750150E+00+1.06143554E-02-3.57999360E-06+5.50363760E-10-3.17051769E-14    2
-6.92747939E+03-1.53833428E+01+2.59479867E+00+2.27100669E-02-1.39473846E-05    3
+4.70095591E-09-6.90044236E-13-4.91486975E+03+1.43240718E+01+0.00000000E+00    4
SC2H4OH    8/12/15      C   2H   5O   1    0G   300.000  5000.000 1385.000     2
+8.15007136E+00+1.02549305E-02-3.40137764E-06+5.17509965E-10-2.96128942E-14    2
-1.05014386E+04-1.73134615E+01+1.46281093E+00+2.39193995E-02-1.30667185E-05    3
+3.10615465E-09-1.85896007E-13-8.00790323E+03+1.92547092E+01+0.00000000E+00    4
O2C2H4OH   9/ 1/12 THERMC   2H   5O   3    0G   300.000  5000.000 1506.000    41
+1.27503881E+01+1.11514325E-02-3.83473891E-06+5.98155829E-10-3.48372108E-14    2
-2.52770876E+04-3.54317608E+01+7.04009800E+00+1.59564166E-02+2.21097416E-06    3
-7.05197355E-09+2.08266026E-12-2.24524432E+04-1.75361758E+00+0.00000000E+00    4
C2H4O2H    9/ 1/12      C   2H   5O   2    0G   300.000  5000.000 1389.000    31
+1.00590614E+01+1.13378955E-02-3.89403387E-06+6.06090687E-10-3.52212353E-14    2
+4.24048653E+02-2.32086536E+01+2.75788364E+00+2.88271987E-02-2.08302264E-05    3
+8.47401397E-09-1.48617610E-12+3.00153893E+03+1.59921711E+01+0.00000000E+00    4
C2H4O1-2          L 8/88C  2 H  4 O  1    0 G   200.000  6000.00  1000.00      1
+5.48876410E+00+1.20461900E-02-4.33369310E-06+7.00283110E-10-4.19490880E-14    2
-9.18042510E+03-7.07996050E+00+3.75905320E+00-9.44121800E-03+8.03097210E-05    3
-1.00807880E-07+4.00399210E-11-7.56081430E+03+7.84974750E+00-6.33046570E+03    4
C2H3O1-2          A 1/05C  2 H  3 O  1    0 G   200.000  6000.00  1000.00      1
+5.60158035E+00+9.17613962E-03-3.28028902E-06+5.27903888E-10-3.15362241E-14    2
+1.71446252E+04-5.47228512E+00+3.58349017E+00-6.02275805E-03+6.32426867E-05    3
-8.18540707E-08+3.30444505E-11+1.85681353E+04+9.59725926E+00+1.97814471E+04    4
CH3CHO            L 8/88C  2 H  4 O   1   0 G   200.000  6000.00  1000.00      1
+5.40411080E+00+1.17230590E-02-4.22631370E-06+6.83724510E-10-4.09848630E-14    2
-2.25931220E+04-3.48079170E+00+4.72945950E+00-3.19328580E-03+4.75349210E-05    3
-5.74586110E-08+2.19311120E-11-2.15728780E+04+4.10301590E+00-1.99879490E+04    4
CH3CO             IU2/03C  2 H  3 O  1    0 G   200.000  6000.00  1000.00      1
+5.31371650E+00+9.17377930E-03-3.32203860E-06+5.39474560E-10-3.24523680E-14    2
-3.64504140E+03-1.67575580E+00+4.03587050E+00+8.77294870E-04+3.07100100E-05    3
-3.92475650E-08+1.52968690E-11-2.68207380E+03+7.86176820E+00-1.23880390E+03    4
CH2CHO            T03/10C  2 H  3 O  1    0 G   200.000  6000.00  1000.00      1
+6.53928338E+00+7.80238629E-03-2.76413612E-06+4.42098906E-10-2.62954290E-14    2
-1.18858659E+03-8.72091393E+00+2.79502600E+00+1.01099472E-02+1.61750645E-05    3
-3.10303145E-08+1.39436139E-11+1.62944975E+02+1.23646657E+01+1.53380440E+03    4
O2CH2CHO          BOZ_03C   2H   3O   3    0G   300.000  5000.000 1393.000    01
+1.11807543E+01+9.14479256E-03-3.15089833E-06+4.91944238E-10-2.86639180E-14    2
-1.55790331E+04-2.87892740E+01-1.29465843E+00+4.44936393E-02-4.26577074E-05    3
+2.07391950E-08-3.96828771E-12-1.18275628E+04+3.60778797E+01+0.00000000E+00    4
HO2CH2CO          BOZ_03C   2H   3O   3    0G   300.000  5000.000 1386.000    01
+1.04146322E+01+1.12680116E-02-5.17494839E-06+1.00333285E-09-6.68165911E-14    2
-1.40955672E+04-2.27894400E+01+2.22681686E+00+3.56781380E-02-3.26401909E-05    3
+1.47651988E-08-2.64794380E-12-1.18735095E+04+1.91581197E+01+0.00000000E+00    4
C2H3OH     2/ 3/ 9 THERMC   2H   4O   1    0G   300.000  5000.000 1410.000    11
+8.32598158E+00+8.03387281E-03-2.63928405E-06+3.98410726E-10-2.26551155E-14    2
-1.83221436E+04-2.02080305E+01-1.27972260E-01+3.38506073E-02-3.30644935E-05    3
+1.64858739E-08-3.19935455E-12-1.59914544E+04+2.30438601E+01+0.00000000E+00    4
C2H2OH                  H   3C   2O   1    0G   300.000  5000.000 1401.000    11
+8.20268447E+00+5.92989165E-03-1.99194448E-06+3.05794341E-10-1.76114732E-14    2
+1.24881328E+04-1.89670436E+01+6.41642616E-01+2.61903633E-02-2.30385370E-05    3
+1.02804704E-08-1.81971416E-12+1.48276951E+04+2.06750999E+01+0.00000000E+00    4
CH2CO     11/13/18 THERMC   2H   2O   1    0G   300.000  5000.000 1400.000     1
 6.32896692E+00 5.44012978E-03-1.82687969E-06 2.80010787E-10-1.60964160E-14    2
-8.36526176E+03-9.53528539E+00 2.35724171E+00 1.62213064E-02-1.34812364E-05    3
 6.11939897E-09-1.13613089E-12-7.11393356E+03 1.12990053E+01                   4
HCCO              T 4/09H  1 C  2 O  1    0 G   200.000  6000.00  1000.00      1
+5.91479333E+00+3.71408730E-03-1.30137010E-06+2.06473345E-10-1.21476759E-14    2
+1.93596301E+04-5.50567269E+00+1.87607969E+00+2.21205418E-02-3.58869325E-05    3
+3.05402541E-08-1.01281069E-11+2.01633840E+04+1.36968290E+01+2.14444387E+04    4
HCCOH             T12/09C  2 H  2 O  1    0 G   200.000  6000.00  1000.00      1
+6.37509678E+00+5.49429011E-03-1.88136576E-06+2.93803536E-10-1.71771901E-14    2
+8.93277676E+03-8.24498007E+00+2.05541154E+00+2.52003372E-02-3.80821654E-05    3
+3.09890632E-08-9.89799902E-12+9.76872113E+03+1.22271534E+01+1.12217316E+04    4
CH3CO3H    6/26/95 THERMC   2H   4O   3    0G   300.000  5000.000 1391.000    31
+1.25060485E+01+9.47789695E-03-3.30402246E-06+5.19630793E-10-3.04233568E-14    2
-4.59856703E+04-3.79195947E+01+2.24135876E+00+3.37963514E-02-2.53887482E-05    3
+9.67583587E-09-1.49266157E-12-4.24677831E+04+1.70668133E+01+0.00000000E+00    4
CH3CO3     4/ 3/ 0 THERMC   2H   3O   3    0G   300.000  5000.000 1391.000    21
+1.12522498E+01+8.33652672E-03-2.89014530E-06+4.52781734E-10-2.64354456E-14    2
-2.60238584E+04-2.96370457E+01+3.60373432E+00+2.70080341E-02-2.08293438E-05    3
+8.50541104E-09-1.43846110E-12-2.34205171E+04+1.12014914E+01+0.00000000E+00    4
CH3CO2     2/14/95 THERMC   2H   3O   2    0G   300.000  5000.000 1395.000    11
+8.54059736E+00+8.32951214E-03-2.84722010E-06+4.41927196E-10-2.56373394E-14    2
-2.97290678E+04-2.03883545E+01+1.37440768E+00+2.49115604E-02-1.74308894E-05    3
+6.24799508E-09-9.09516835E-13-2.72330150E+04+1.81405454E+01+0.00000000E+00    4
CH3OCH3                 H  6 C  2 O  1      G     298.0    3000.0    1000.0    1
+1.13851970E+00+2.58202899E-02-1.29425822E-05+3.14818537E-09-3.01294764E-13    2
-2.35157473E+04+1.85133202E+01+3.75480003E+00+9.94330522E-03+2.04658920E-05    3
-2.65048607E-08+9.20398140E-12-2.38174871E+04+7.12147313E+00+0.00000000E+00    4
CH3OCH2                 H  5 C  2 O  1      G     298.0    3000.0    1000.0    1
+2.74300130E+00+2.06529566E-02-1.03925669E-05+2.54086134E-09-2.44516053E-13    2
-1.32986515E+03+1.24007048E+01+3.93734319E+00+9.90763869E-03+1.63345997E-05    3
-2.34568933E-08+8.57704791E-12-1.32547779E+03+7.99274498E+00+0.00000000E+00    4
CH3OCH2O2H 2/12/14 THERMC   2H   6O   3    0G   300.000  5000.000 1404.000    31
+1.28159161E+01+1.34818095E-02-4.50397729E-06+6.88229286E-10-3.94883680E-14    2
-4.06745921E+04-3.78047802E+01+1.05786981E+00+4.36787095E-02-3.46383899E-05    3
+1.44808830E-08-2.46100643E-12-3.68851076E+04+2.43391936E+01+0.00000000E+00    4
CH3OCH2O2  2/12/14 THERMC   2H   5O   3    0G   300.000  5000.000 1441.000    21
+1.19179361E+01+1.19412867E-02-3.93526185E-06+5.95756132E-10-3.39597705E-14    2
-2.34231833E+04-3.20096863E+01+3.39930541E+00+3.09460407E-02-1.92548181E-05    3
+5.76033887E-09-6.16081571E-13-2.04433218E+04+1.39429608E+01+0.00000000E+00    4
CH2OCH2O2H 2/12/14 THERMC   2H   5O   3    0G   300.000  5000.000 1418.000    21
+1.23892901E+01+1.11758961E-02-3.59249095E-06+5.34196366E-10-3.00536541E-14    2
-1.80551598E+04-3.29576862E+01+1.62245477E-01+4.76101093E-02-4.52046954E-05    3
+2.18379311E-08-4.11295947E-12-1.46498100E+04+2.98253164E+01+0.00000000E+00    4
O2CH2OCH2O2H 2/12/14 ERMC   2H   5O   5    0G   300.000  5000.000 1433.000    31
+1.77378326E+01+1.13589899E-02-3.67382539E-06+5.49255712E-10-3.10405899E-14    2
-3.82903058E+04-5.66609932E+01+2.39977678E+00+5.39881943E-02-4.87969524E-05    3
+2.19792134E-08-3.86106979E-12-3.37824638E+04+2.30683371E+01+0.00000000E+00    4
HO2CH2OCHO 2/12/14 THERMC   2H   4O   4    0G   300.000  5000.000 1386.000    31
+1.57136128E+01+9.64430166E-03-3.44136025E-06+5.49722196E-10-3.25360322E-14    2
-6.29409094E+04-5.29505242E+01+1.21909586E+00+4.28858235E-02-3.17634222E-05    3
+1.11542676E-08-1.49753153E-12-5.79287926E+04+2.49759193E+01+0.00000000E+00    4
OCH2OCHO   5/29/14 THERMC   2H   3O   3    0G   300.000  5000.000 1523.000    21
+1.24013200E+01+7.83738243E-03-2.82992688E-06+4.55558739E-10-2.71061389E-14    2
-4.68453470E+04-3.78084549E+01+1.89539692E+00+2.74118545E-02-1.36476090E-05    3
+1.26325603E-09+5.17970476E-13-4.27879440E+04+2.02333278E+01+0.00000000E+00    4
HOCH2OCO   5/29/14 THERMC   2H   3O   3    0G   300.000  5000.000 1443.000    11
+1.11498410E+01+9.34736520E-03-3.35541548E-06+5.38037115E-10-3.19260183E-14    2
-4.75012119E+04-2.95983867E+01+5.95255071E+00+8.42196282E-03+1.36741678E-05    3
-1.46786275E-08+3.84143533E-12-4.44470269E+04+2.85657217E+00+0.00000000E+00    4
CH3OCH2OH  2/ 9/96 THERMC   2H   6O   2    0G   300.000  5000.000 2014.000    31
+8.70981570E+00+1.53602372E-02-5.41003788E-06+8.60573446E-10-5.08819752E-14    2
-4.76607115E+04-1.80226702E+01+3.15851876E+00+2.44325751E-02-8.66984784E-06    3
-5.93319328E-11+4.36400003E-13-4.54488899E+04+1.30511235E+01+0.00000000E+00    4
CH3OCH2O   5/15/14 THERMC   2H   5O   2    0G   300.000  5000.000 1523.000    31
+9.81288609E+00+1.21313106E-02-4.30285768E-06+6.84443177E-10-4.03862658E-14    2
-2.50760742E+04-2.51866352E+01+5.63414373E+00+8.92830283E-03+1.37225633E-05    3
-1.40497059E-08+3.54625624E-12-2.22825214E+04+1.93588846E+00+0.00000000E+00    4
CH3OCHO                 H  4 C  2 O  2      G     298.0    3000.0    1000.0    1 !\AUTHOR: KPS !\REF: DAMES, CNF, 2016 !\COMMENT:
+1.55821560E+00+2.63651102E-02-1.49021985E-05+3.93577994E-09-3.99334221E-13    2
-4.47996443E+04+1.82846496E+01+3.95242735E+00+6.27936769E-03+3.21013314E-05    3
-3.93941104E-08+1.36185570E-11-4.47899337E+04+9.26882234E+00+0.00000000E+00    4
CH3OCO                  H  3 C  2 O  2      G     298.0    3000.0    1000.0    1 !\AUTHOR: KPS !\REF: DAMES, CNF, 2016 !\COMMENT:
+3.36304128E+00+1.87670995E-02-1.03048118E-05+2.67955225E-09-2.69524760E-13    2
-2.08317053E+04+1.09017923E+01+4.20427121E+00+8.77414983E-03+1.52020481E-05    3
-2.17223880E-08+7.77727542E-12-2.06876220E+04+8.45258172E+00+0.00000000E+00    4
CH2OCHO                 H  3 C  2 O  2      G     298.0    3000.0    1000.0    1 !\AUTHOR: KPS !\REF: DAMES, CNF, 2016 !\COMMENT:
+5.66297823E+00+1.73979570E-02-1.01218468E-05+2.73226211E-09-2.81907442E-13    2
-2.14389479E+04-2.38514196E+00+3.19932230E+00+1.93736375E-02-1.21521306E-06    3
-1.11559169E-08+5.18761324E-12-2.05538696E+04+1.14662057E+01+0.00000000E+00    4
C3H8       8/12/15      C   3H   8    0    0G   300.000  5000.000 1390.000    21
+9.15541310E+00+1.72574139E-02-5.85614868E-06+9.04190155E-10-5.22523772E-14    2
-1.75762439E+04-2.77418510E+01+2.40878470E-01+3.39548599E-02-1.60930874E-05    3
+2.83480628E-09+2.78195172E-14-1.40362853E+04+2.16500800E+01+0.00000000E+00    4
IC3H7      8/12/15      C   3H   7    0    0G     298.0    6000.0    1000.0    1
+6.70775549E+00+1.74048076E-02-6.07615926E-06+9.60084351E-10-5.65656490E-14    2
+7.55377821E+03-1.03686516E+01-8.97467137E-01+4.15744022E-02-4.94778349E-05    3
+4.56493655E-08-1.79085437E-11+9.93950407E+03+2.92641758E+01+0.00000000E+00    4
NC3H7      8/12/15      C   3H   7    0    0G     298.0    6000.0    1000.0    1
+7.48614243E+00+1.65769478E-02-5.74876481E-06+9.04103694E-10-5.30867231E-14    2
+8.93710008E+03-1.42595379E+01-2.20120865E+00+5.29641653E-02-7.23640506E-05    3
+6.36996940E-08-2.29332581E-11+1.15130744E+04+3.43669174E+01+0.00000000E+00    4
NC3H7O2H   8/12/15      C   3H   8O   2    0G   300.000  5000.000 1392.000    41
+1.42246236E+01+1.74340964E-02-5.97063522E-06+9.27753851E-10-5.38585168E-14    2
-2.88159737E+04-4.74357865E+01+1.35815897E+00+4.56683952E-02-2.91646368E-05    3
+9.41701313E-09-1.22337394E-12-2.41528416E+04+2.23322825E+01+0.00000000E+00    4
NC3H7O2    8/12/15      C   3H   7O   2    0G   300.000  5000.000 1390.000    31
+1.32753283E+01+1.61303126E-02-5.52348308E-06+8.58197168E-10-4.98172586E-14    2
-1.16032968E+04-4.15091215E+01+2.13311681E+00+3.96692045E-02-2.37570127E-05    3
+6.96020417E-09-7.82576856E-13-7.46687112E+03+1.92444565E+01+0.00000000E+00    4
IC3H7O2H   8/12/15      C   3H   8O   2    0G   300.000  5000.000 1405.000    41
+1.44896107E+01+1.68268026E-02-5.67601391E-06+8.72850837E-10-5.02993991E-14    2
-3.06478491E+04-5.01352281E+01+1.77384705E+00+4.75813498E-02-3.43745304E-05    3
+1.31405381E-08-2.06922904E-12-2.63458844E+04+1.77669753E+01+0.00000000E+00    4
IC3H7O2    8/12/15      C   3H   7O   2    0G   300.000  5000.000 1407.000    31
+1.35268120E+01+1.54306581E-02-5.17464218E-06+7.92548669E-10-4.55415379E-14    2
-1.33946348E+04-4.40461451E+01+2.58517502E+00+4.16107259E-02-2.92193877E-05    3
+1.08614807E-08-1.66312005E-12-9.67013161E+03+1.44731300E+01+0.00000000E+00    4
C3H6OOH1-2 9/ 1/12      C   3H   7O   2    0G   300.000  5000.000 1387.000    41
+1.38088686E+01+1.43845650E-02-4.74440961E-06+7.19308280E-10-4.10654123E-14    2
-5.14352831E+03-4.20210765E+01+2.83631132E+00+3.88229894E-02-2.47944364E-05    3
+7.85644898E-09-9.58634300E-13-1.26002528E+03+1.72549973E+01+0.00000000E+00    4
C3H6OOH1-3 9/ 1/12      C   3H   7O   2    0G   300.000  5000.000 1401.000    41
+1.39130757E+01+1.40218463E-02-4.55921149E-06+6.84182417E-10-3.87696213E-14    2
-3.65650518E+03-4.21532559E+01+1.74271107E+00+4.53733504E-02-3.57580373E-05    3
+1.48540053E-08-2.49981756E-12+2.32580844E+02+2.20973041E+01+0.00000000E+00    4
C3H6OOH2-1 9/ 1/12      C   3H   7O   2    0G   300.000  5000.000 1393.000    41
+1.36645362E+01+1.54329764E-02-5.29285952E-06+8.23001262E-10-4.77931121E-14    2
-5.58295862E+03-4.28758364E+01+2.38465746E+00+4.42928555E-02-3.50977087E-05    3
+1.53695144E-08-2.81167824E-12-1.80979612E+03+1.69923285E+01+0.00000000E+00    4
C3H6OOH1-2O2 9/ 1/12    C   3H   7O   4    0G   300.000  5000.000 1404.000    51
+1.91044980E+01+1.44076100E-02-4.72127814E-06+7.12631642E-10-4.05578490E-14    2
-2.50270510E+04-6.63747978E+01+3.99085043E+00+5.31865338E-02-4.28597948E-05    3
+1.77187019E-08-2.92768695E-12-2.02143526E+04+1.34150719E+01+0.00000000E+00    4
C3H6OOH1-3O2 9/ 1/12    C   3H   7O   4    0G   300.000  5000.000 1416.000    51
+1.81661664E+01+1.47644887E-02-4.74842743E-06+7.06972467E-10-3.98305587E-14    2
-2.26256376E+04-5.93719393E+01+5.56933350E+00+4.68523421E-02-3.58917784E-05    3
+1.43314525E-08-2.29776083E-12-1.86065694E+04+7.18655005E+00+0.00000000E+00    4
C3H6OOH2-1O2 9/ 1/12    C   3H   7O   4    0G   300.000  5000.000 1404.000    51
+1.91044980E+01+1.44076100E-02-4.72127814E-06+7.12631642E-10-4.05578490E-14    2
-2.50270510E+04-6.63747978E+01+3.99085043E+00+5.31865338E-02-4.28597948E-05    3
+1.77187019E-08-2.92768695E-12-2.02143526E+04+1.34150719E+01+0.00000000E+00    4
C3H5-1E-2OOH            C  3 H  6 O  2      G     298.0    6000.0    1000.0    1
 1.25352860E+01 1.41801036E-02-4.86408170E-06 7.59244931E-10-4.43443519E-14    2
-1.42746980E+04-3.75622448E+01-1.92214080E+00 7.47575190E-02-1.14477005E-04    3
 9.60658373E-08-3.18580028E-11-1.10322543E+04 3.27197181E+01                   4
C3KET12   10/17/12      C   3H   6O   3    0G   300.000  5000.000 1385.000    41
+1.70187760E+01+1.32097361E-02-4.67054741E-06+7.41411770E-10-4.36869787E-14    2
-4.23572589E+04-5.92615939E+01+1.03882879E+00+5.34180080E-02-4.47684141E-05    3
+1.94651680E-08-3.45055244E-12-3.70308881E+04+2.56511209E+01+0.00000000E+00    4
C3KET13   10/17/12      C   3H   6O   3    0G   300.000  5000.000 1508.000    41
+1.73612692E+01+1.32330813E-02-4.75332110E-06+7.62529227E-10-4.52613717E-14    2
-4.06248060E+04-6.17768199E+01+4.74956819E+00+3.14080991E-02-6.83838427E-06    3
-5.67123901E-09+2.27686972E-12-3.51924570E+04+9.83753744E+00+0.00000000E+00    4
C3H51-2,3OOH 8/26/3 THRMC   3H   7O   4    0G   300.000  5000.000 1386.000    61
+2.12378169E+01+1.39519596E-02-4.94539222E-06+7.86381389E-10-4.63925564E-14    2
-1.92864584E+04-7.69636561E+01+2.55619708E+00+6.13504487E-02-5.23205391E-05    3
+2.28208029E-08-4.02231508E-12-1.31353414E+04+2.21043799E+01+0.00000000E+00    4
C3H52-1,3OOH 8/26/3 THRMC   3H   7O   4    0G   300.000  5000.000 1379.000    61
+2.02817964E+01+1.48155431E-02-5.25503386E-06+8.35963453E-10-4.93308915E-14    2
-1.80085066E+04-7.22688262E+01+4.12253742E+00+5.19553611E-02-3.83733727E-05    3
+1.45851637E-08-2.29820536E-12-1.22759164E+04+1.48367359E+01+0.00000000E+00    4
C3H5O1-2OOH-3 10/13 THERC   3H   6O   3    0G   300.000  5000.000 1432.000    31
+1.57042382E+01+1.30255692E-02-4.23544254E-06+6.35555595E-10-3.60110207E-14    2
-2.77269333E+04-5.51895464E+01-3.25001215E+00+6.65787151E-02-6.18859778E-05    3
+2.84638649E-08-5.08511634E-12-2.22371240E+04+4.30381280E+01+0.00000000E+00    4
C3H5O1-3OOH-2 10/13 THERC   3H   6O   3    0G   300.000  5000.000 1434.000    21
+1.44493479E+01+1.36372560E-02-4.25836513E-06+6.20006211E-10-3.43451580E-14    2
-2.77372360E+04-5.06099103E+01-4.43959178E+00+7.16532928E-02-7.15032351E-05    3
+3.51737842E-08-6.63682938E-12-2.27250412E+04+4.56394038E+01+0.00000000E+00    4
C3H6O1-2          A01/05C  3 H  6 O  1    0 G   200.000  6000.00  1000.00      1
+8.01491079E+00+1.73919953E-02-6.26027968E-06+1.01188256E-09-6.06239111E-14    2
-1.51980838E+04-1.88279964E+01+3.42806676E+00+6.25176642E-03+6.13196311E-05    3
-8.60387185E-08+3.51371393E-11-1.28446646E+04+1.04244994E+01-1.11564001E+04    4
C3H6O1-3          A11/04C  3 H  6 O  1    0 G   200.000  6000.00  1000.00      1
+6.80716906E+00+1.88824545E-02-6.79082475E-06+1.09713919E-09-6.57154952E-14    2
-1.36547629E+04-1.35382154E+01+5.15283752E+00-1.86401716E-02+1.29980652E-04    3
-1.58629974E-07+6.20668783E-11-1.13243512E+04+4.73561224E+00-9.75233898E+03    4
C3H5-SOOH               C  3 H  6 O  2      G     298.0    6000.0    1000.0    1
 1.17366777E+01 1.50781115E-02-5.22873766E-06 8.22569776E-10-4.83198810E-14    2
-1.19051570E+04-3.21649975E+01 6.05480242E-03 5.72962550E-02-7.65094431E-05    3
 6.36300985E-08-2.20626642E-11-8.82238404E+03 2.68572270E+01                   4
C3H6       8/12/15      C   3H   6    0    0G   298.000  6000.000 1000.000    01
+6.59032304E+00+1.52592866E-02-5.30369441E-06+8.35510888E-10-4.91215549E-14    2
-2.47481113E+02-1.15748238E+01-1.54606737E+00+4.36553128E-02-5.61392417E-05    3
+4.98421927E-08-1.84798923E-11+2.07056233E+03+2.99232495E+01+0.00000000E+00    4
C3H5-A     8/12/15      C   3H   5    0    0G   298.000  6000.000 1000.000    01
+7.37604097E+00+1.23449782E-02-4.26463882E-06+6.69045835E-10-3.92202554E-14    2
+1.77332960E+04-1.61758204E+01-3.32899442E+00+5.38423469E-02-7.65500752E-05    3
+6.35512285E-08-2.14283003E-11+2.03420628E+04+3.68038362E+01+0.00000000E+00    4
C3H5-S     8/12/15      C   3H   5    0    0G   300.000  5000.000 1390.000    11
+7.95954498E+00+1.11163183E-02-3.75197834E-06+5.77246260E-10-3.32768957E-14    2
+2.80567891E+04-1.79800372E+01+1.61793372E+00+2.44803904E-02-1.41856503E-05    3
+4.16402233E-09-4.90904795E-13+3.04291037E+04+1.66341443E+01+0.00000000E+00    4
C3H5-T     8/12/15      C   3H   5    0    0G   300.000  5000.000 1376.000    11
+7.69949212E+00+1.17803985E-02-4.07791749E-06+6.38119222E-10-3.72229675E-14    2
+2.61747145E+04-1.68305890E+01+2.29256998E+00+1.98527646E-02-6.42635654E-06    3
-5.90016395E-10+5.05491095E-13+2.85773377E+04+1.39407124E+01+0.00000000E+00    4
CC3H6                   C   3H   6O   0    0G   200.000  6000.000 1000.        1
+6.21663437E+00+1.65393591E-02-5.90075838E-06+9.48095199E-10-5.65661522E-14    2
+2.95937491E+03-1.36041009E+01+2.83278674E+00-5.21028618E-03+9.29583210E-05    3
-1.22753194E-07+4.99191366E-11+5.19520048E+03+1.08306333E+01+6.41047999E+03    4
CH3CHCHO                C   3H   5O   1    0G   300.000  5000.000 1424.000    21
+1.06781476E+01+1.12805711E-02-3.89010759E-06+6.07617268E-10-3.54120848E-14    2
-7.73234209E+03-3.24971238E+01+1.47166733E+00+2.69251618E-02-1.00248013E-05    3
-1.13421435E-09+1.03416658E-12-4.04142023E+03+1.88722472E+01+0.00000000E+00    4
CH3CHCO   03/03/95 THERMC   3H   4O   1    0G   300.000  5000.000 1400.00     41
+1.00219123E+01+9.56966300E-03-3.26221644E-06+5.05231706E-10-2.92593257E-14    2
-1.42482738E+04-2.77829973E+01+1.48380119E+00+3.22203013E-02-2.70250033E-05    3
+1.20499164E-08-2.18365931E-12-1.15276540E+04+1.71552068E+01+0.00000000E+00    4
C3H5O             KPS12 C   3H   5O   1    0G   300.000  5000.000 1402.000    01
+1.02638186E+01+1.17609932E-02-3.89837957E-06+5.92650815E-10-3.38867417E-14    2
+7.25938472E+03-2.75108651E+01+8.24068673E-01+3.46749909E-02-2.51786795E-05    3
+9.56781953E-09-1.48085302E-12+1.04203725E+04+2.28283070E+01+0.00000000E+00    4
CH2CHOCH2  8/ 8/15      C   3H   5O   1    0G   300.000  5000.000 1384.000    21
+1.20076931E+01+1.05055204E-02-3.69920541E-06+5.85629983E-10-3.44431587E-14    2
+6.97311613E+03-3.75189859E+01+1.15350351E+00+3.51253596E-02-2.50071619E-05    3
+9.00715632E-09-1.32376643E-12+1.08300872E+04+2.10606652E+01+0.00000000E+00    4
AC4H7OOH   6/17/13 THERMC   4H   8O   2    0G   300.000  5000.000 1395.000    41
+1.47661443E+01+2.12235231E-02-7.09403390E-06+1.08423759E-09-6.22145708E-14    2
-1.35617411E+04-4.77449138E+01+1.33470633E+00+5.27831440E-02-3.58861360E-05    3
+1.32495013E-08-2.06619289E-12-8.87891782E+03+2.43857336E+01+0.00000000E+00    4
AC3H5OOH    GOLDSMITH   C   3H   6O   2    0G   298.0    6000.0   1000.000    31
+1.20838649E+01+1.47946591E-02-5.13212591E-06+8.07504999E-10-4.74394983E-14    2
-1.02184463E+04-3.36434791E+01+3.18124993E+00+4.35233041E-02-5.16277353E-05    3
+4.32011427E-08-1.57714983E-11-7.63521503E+03+1.21725683E+01+0.00000000E+00    4
C3H4-P            T 2/90H  4 C  3    0    0 G   200.000  6000.00  1000.00      1
+6.02524000E+00+1.13365420E-02-4.02233910E-06+6.43760630E-10-3.82996350E-14    2
+1.96209420E+04-8.60437850E+00+2.68038690E+00+1.57996510E-02+2.50705960E-06    3
-1.36576230E-08+6.61542850E-12+2.08023740E+04+9.87693510E+00+2.23020590E+04    4
C3H4-A            L 8/89C  3 H  4    0    0 G   200.000  6000.00  1000.00      1
+6.31687220E+00+1.11337280E-02-3.96293780E-06+6.35642380E-10-3.78755400E-14    2
+2.01174950E+04-1.09957660E+01+2.61304450E+00+1.21225750E-02+1.85398800E-05    3
-3.45251490E-08+1.53350790E-11+2.15415670E+04+1.02261390E+01+2.29622670E+04    4
C3H3              T 7/11C  3 H  3    0    0 G   200.000  6000.00  1000.000     1
+7.14221719E+00+7.61902211E-03-2.67460030E-06+4.24914904E-10-2.51475443E-14    2
+3.95709594E+04-1.25848690E+01+1.35110873E+00+3.27411291E-02-4.73827407E-05    3
+3.76310220E-08-1.18541128E-11+4.07679941E+04+1.52058598E+01+4.22762135E+04    4
CC3H4             T12/81C   3H   4    0    0G   300.000  5000.00  1000.00      1
+6.69999310E+00+1.03573720E-02-3.45511670E-06+5.06529490E-10-2.66822760E-14    2
+3.01990510E+04-1.33787700E+01-2.46210470E-02+2.31972150E-02-1.84743570E-06    3
-1.59275930E-08+8.68461550E-12+3.23341370E+04+2.27297620E+01+3.33272800E+04    4
C3H2              T12/00C  3 H  2    0    0 G   200.000  6000.00  1000.00      1
+6.67324762E+00+5.57728845E-03-1.99180164E-06+3.20289156E-10-1.91216272E-14    2
+7.57571184E+04-9.72894405E+00+2.43417332E+00+1.73013063E-02-1.18294047E-05    3
+1.02756396E-09+1.62626314E-12+7.69074892E+04+1.21012230E+01+7.83005132E+04    4
H2CCC(S)               0C   3H   2    0    0G   200.000  5000.000 1500.00    0 1
+6.48887620E+00+5.31127890E-03-1.78094900E-06+2.72526420E-10-1.56195900E-14    2
+6.36618640E+04-1.00642830E+01+3.72297260E+00+9.25898540E-03-2.30061910E-06    3
-1.02008080E-09+4.53743570E-13+6.48772890E+04+5.68659360E+00+0.00000000E+00    4
C3H2(S)                0C   3H   2    0    0G   200.000  5000.000  900.00    0 1
+7.76425700E+00+4.71127740E-03-1.61706370E-06+2.54724060E-10-1.50385720E-14    2
+6.68496720E+04-1.50985490E+01+5.29764820E+00+1.69874660E-02-2.42665170E-05    3
+1.86536810E-08-5.57630010E-12+6.72404660E+04-3.75400410E+00+0.00000000E+00    4
C3H2C                  0C   3H   2    0    0G   200.000  5000.000 1500.00    0 1
+6.56326800E+00+5.23632560E-03-1.75448300E-06+2.68661060E-10-1.54285090E-14    2
+5.65146180E+04-1.20006070E+01+1.12958880E+00+1.72874010E-02-1.13668230E-05    3
+3.45692960E-09-3.66159510E-13+5.84190800E+04+1.73314480E+01+0.00000000E+00    4
PC3H4OH-1  9/25/15      C   3H   5O   1    0G   300.000  5000.000 1403.000    21
+1.09468986E+01+1.04014540E-02-3.44082448E-06+5.22105632E-10-2.98049266E-14    2
+4.11530600E+03-3.11161699E+01+2.07150195E+00+3.50016810E-02-3.01922013E-05    3
+1.38467853E-08-2.55380109E-12+6.81914209E+03+1.51916605E+01+0.00000000E+00    4
PC3H4OH-2  4/ 2/13 THERMC   3H   5O   1    0G   300.000  5000.000 1403.000    21
+1.07164095E+01+1.06066461E-02-3.51374060E-06+5.33713932E-10-3.04901511E-14    2
+4.98486803E+03-2.98329329E+01+1.42757363E+00+3.64825569E-02-3.18007132E-05    3
+1.46914605E-08-2.72331227E-12+7.80342663E+03+1.85890339E+01+0.00000000E+00    4
PC3H4OH-3  9/25/15      C   3H   5O   1    0G   300.000  5000.000 1378.000    11
+1.15297558E+01+1.14381097E-02-4.04415495E-06+6.41949269E-10-3.78242456E-14    2
-3.45486444E+03-3.65385497E+01+4.06368169E-01+3.70231405E-02-2.72202689E-05    3
+1.05783475E-08-1.73632514E-12+5.27160824E+02+2.34781848E+01+0.00000000E+00    4
SC3H4OH    3/28/13      C   3H   5O   1    0G   300.000  5000.000 1407.000    21
+1.20968484E+01+9.43976596E-03-3.10773897E-06+4.69609188E-10-2.67165710E-14    2
-3.85854894E+02-3.76795997E+01+1.72870561E+00+4.41015870E-02-4.72013860E-05    3
+2.52073596E-08-5.13375710E-12+2.22720503E+03+1.43928257E+01+0.00000000E+00    4
C3H3O      2/17/14 CZHOUH   3C   3O   1     G   298.150  2000.000 1000.00      1
+4.19355696E+00+1.95625103E-02-1.22336450E-05+3.90615061E-09-5.08539231E-13    2
+3.14931737E+04+5.03216224E+00+8.75023836E-01+3.51184068E-02-3.89901356E-05    3
+2.40255750E-08-6.10883631E-12+3.20427921E+04+2.04717253E+01+0.00000000E+00    4
C3H3O2H    1/31/13      C   3H   4O   2    0G   300.000  5000.000 1385.000    31
+1.38152174E+01+8.62174763E-03-3.06710006E-06+4.88874247E-10-2.88888385E-14    2
+6.29182941E+03-4.39151257E+01+1.09787313E+00+4.22717882E-02-3.83969355E-05    3
+1.77405069E-08-3.27674312E-12+1.03592314E+04+2.30651783E+01+0.00000000E+00    4
C2HCHO     1/31/13      C   3H   2O   1    0G   300.000  5000.000 2012.000    11
+7.99952054E+00+7.07825497E-03-2.63086819E-06+4.33073185E-10-2.62003284E-14    2
+8.71863156E+03-1.57226237E+01+4.20776611E+00+1.34382727E-02-5.15442099E-06    3
-2.24570818E-11+2.74111284E-13+1.02117375E+04+5.43871873E+00+0.00000000E+00    4
NC3H7OH    3/22/16 THERMC   3H   8O   1    0G   300.000  5000.000 1403.000    11 ! PAWEL ADDED PROPONAL 27/06/2016 
+1.12833724E+01+1.71531932E-02-5.56084500E-06+8.32706677E-10-4.71118622E-14    2
-3.64174301E+04-3.37180466E+01+5.70007484E-02+4.17375704E-02-2.49234034E-05    3
+7.16029301E-09-7.25069606E-13-3.24306821E+04+2.70290017E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 27/06/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 27/06/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1 10/ 2/15      C   3H   7O   1    0G   300.000  5000.000 1388.000    31
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 11/03/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1 10/ 2/15      C   3H   7O   1    0G   300.000  5000.000 1388.000    31
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 11/03/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 27/06/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 27/06/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1 10/ 2/15      C   3H   7O   1    0G   300.000  5000.000 1388.000    31
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 11/03/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1 10/ 2/15      C   3H   7O   1    0G   300.000  5000.000 1388.000    31
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 11/03/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 27/06/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 27/06/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1 10/ 2/15      C   3H   7O   1    0G   300.000  5000.000 1388.000    31
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 11/03/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1 10/ 2/15      C   3H   7O   1    0G   300.000  5000.000 1388.000    31
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 11/03/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 27/06/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 27/06/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1 10/ 2/15      C   3H   7O   1    0G   300.000  5000.000 1388.000    31
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 11/03/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1 10/ 2/15      C   3H   7O   1    0G   300.000  5000.000 1388.000    31
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 11/03/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 27/06/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 27/06/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1 10/ 2/15      C   3H   7O   1    0G   300.000  5000.000 1388.000    31
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 11/03/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1 10/ 2/15      C   3H   7O   1    0G   300.000  5000.000 1388.000    31
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 11/03/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 27/06/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 27/06/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1 10/ 2/15      C   3H   7O   1    0G   300.000  5000.000 1388.000    31
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 11/03/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1 10/ 2/15      C   3H   7O   1    0G   300.000  5000.000 1388.000    31
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 11/03/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 27/06/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 27/06/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1 10/ 2/15      C   3H   7O   1    0G   300.000  5000.000 1388.000    31
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 11/03/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1 10/ 2/15      C   3H   7O   1    0G   300.000  5000.000 1388.000    31
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 11/03/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 27/06/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 27/06/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1 10/ 2/15      C   3H   7O   1    0G   300.000  5000.000 1388.000    31
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 11/03/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1 10/ 2/15      C   3H   7O   1    0G   300.000  5000.000 1388.000    31
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-1  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1388.000    31 ! PAWEL ADDED PROPONAL 11/03/2016 
+1.14795375E+01+1.45881429E-02-4.88359380E-06+7.47606975E-10-4.29608360E-14    2
-1.46832088E+04-3.36825807E+01+1.13614529E+00+3.68850655E-02-2.24073579E-05    3
+6.62398992E-09-7.32206246E-13-1.09273174E+04+2.24919343E+01+0.00000000E+00    4
C3H6OH1-2  9/ 1/12      C   3H   7O   1    0G   300.000  5000.000 1395.000    31
+1.00338281E+01+1.60227373E-02-5.41658448E-06+8.34191172E-10-4.81215988E-14    2
-1.27912397E+04-2.39034395E+01+5.05207596E-01+3.63869988E-02-2.15530901E-05    3
+6.45584786E-09-7.71267046E-13-9.26980840E+03+2.79804349E+01+0.00000000E+00    4
C3H6OH1-3  3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1398.000    31 ! PAWEL ADDED PROPONAL 27/06/2016 
+1.12537269E+01+1.48842686E-02-5.00124819E-06+7.67003856E-10-4.41140957E-14    2
-1.10522005E+04-3.16714219E+01+2.53522975E+00+3.42021055E-02-2.11910432E-05    3
+6.89184707E-09-9.29272171E-13-7.89969902E+03+1.55562988E+01+0.00000000E+00    4
NC3H7O     8/12/15      C   3H   7O   1    0G   300.000  5000.000 1386.000    21
+1.15279177E+01+1.53775991E-02-5.23946272E-06+8.11382512E-10-4.69927603E-14    2
-9.85099867E+03-3.54233008E+01+2.57486880E+00+3.07100600E-02-1.20048836E-05    3
+3.40807108E-12+7.25275283E-13-6.20913350E+03+1.45966401E+01+0.00000000E+00    4
NC3H7O     3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1373.000    31 ! PAWEL ADDED PROPONAL 27/06/2016
+1.20474234E+01+1.49751431E-02-5.20322995E-06+8.16418111E-10-4.77188024E-14    2
-1.01623631E+04-3.85989654E+01+2.49889328E+00+3.08482157E-02-1.17519191E-05    3
-2.91153414E-10+7.87069067E-13-6.19430400E+03+1.49795637E+01+0.00000000E+00    4
C3H5OH            T06/10C  3 H  6 O  1    0 G   200.000  6000.00  1000.00      1
+8.72477114E+00+1.63942712E-02-5.90852993E-06+9.53262253E-10-5.70318010E-14    2
-1.90496618E+04-1.97198674E+01+3.15011905E+00+1.28538274E-02+4.28438434E-05    3
-6.67818707E-08+2.80408237E-11-1.66413668E+04+1.35066359E+01-1.48710589E+04    4
SC3H5OH    2/ 3/ 9      C   3H   6O   1    0G   300.000  5000.000 1404.000    21
+1.11222064E+01+1.27745410E-02-4.25315532E-06+6.48216484E-10-3.71190850E-14    2
-2.36690795E+04-3.41335182E+01-3.53977226E-02+4.34969453E-02-3.74479918E-05    3
+1.70906074E-08-3.13775054E-12-2.02502608E+04+2.41528201E+01+0.00000000E+00    4
CH2CCH2OH  9/ 8/95 THERMC   3H   5O   1    0G   300.000  5000.000 1372.00     21
+9.70702027E+00+1.13972660E-02-3.77993962E-06+5.75209277E-10-3.29229125E-14    2
+9.13212884E+03-2.25012933E+01+2.88422544E+00+2.42428071E-02-1.14152268E-05    3
+1.71775334E-09+1.42177454E-13+1.17935615E+04+1.52102335E+01+0.00000000E+00    4
HOC3H6O2   9/ 1/12      C   3H   7O   3    0G   300.000  5000.000 1407.000    41
+1.56948113E+01+1.57703692E-02-5.30501726E-06+8.14307835E-10-4.68666193E-14    2
-3.24540840E+04-5.06084117E+01+2.84960487E+00+4.77244552E-02-3.60392974E-05    3
+1.43479922E-08-2.33507634E-12-2.82106103E+04+1.76478537E+01+0.00000000E+00    4
IC3H7OH    3/22/16 THERMC   3H   8O   1    0G   300.000  5000.000 1386.000    21 ! PAWEL ADDED PROPONAL 27/06/2016 
+1.25041367E+01+1.62138229E-02-5.35019502E-06+8.11483646E-10-4.63435081E-14    2
-3.89975520E+04-4.25158566E+01+2.53082165E-01+4.17885514E-02-2.38155431E-05    3
+5.85131023E-09-3.55868677E-13-3.45269684E+04+2.42125060E+01+0.00000000E+00    4
C3H6OH2-1  8/ 9/ 4 THERMC   3H   7O   1    0G   300.000  5000.000 1392.000    31
+1.12222277E+01+1.36444398E-02-4.51406709E-06+7.10523275E-10-4.22690392E-14    2
-1.75350136E+04-3.18911926E+01+1.09670360E+00+3.80727565E-02-2.75022497E-05    3
+1.07477493E-08-1.74895773E-12-1.40764487E+04+2.22475799E+01+0.00000000E+00    4
TC3H6OH    8/ 9/ 4 THERMC   3H   7O   1    0G   300.000  5000.000 1392.000    31
+1.12222277E+01+1.36444398E-02-4.51406709E-06+7.10523275E-10-4.22690392E-14    2
-1.75350136E+04-3.18911926E+01+1.09670360E+00+3.80727565E-02-2.75022497E-05    3
+1.07477493E-08-1.74895773E-12-1.40764487E+04+2.22475799E+01+0.00000000E+00    4
TC3H6OH    3/22/16 THERMC   3H   7O   1    0G   300.000  5000.000 1395.000    21 ! PAWEL ADDED PROPONAL 27/06/2016 
+1.11459258E+01+1.48039838E-02-4.85169467E-06+7.31732890E-10-4.16009558E-14    2
-1.67131356E+04-3.26731509E+01+2.20099551E+00+3.52032645E-02-2.24264295E-05    3
+7.53741947E-09-1.04152802E-12-1.35671134E+04+1.55256038E+01+0.00000000E+00    4
IC3H7O     8/12/15      C   3H   7O   1    0G   300.000  5000.000 1527.000    21
+1.19648494E+01+1.42943974E-02-4.71413211E-06+7.14027066E-10-4.07161162E-14    2
-1.17519389E+04-3.88860959E+01+2.36108410E+00+3.45650027E-02-1.94579631E-05    3
+4.71536901E-09-2.64704937E-13-8.28791395E+03+1.33112436E+01+0.00000000E+00    4
IC3H5OH    8/ 1/95 THERMC   3H   6O   1    0G   300.000  5000.000 1374.00     21
+1.07381025E+01+1.31698194E-02-4.41529622E-06+6.77009837E-10-3.89608901E-14    2
-2.47298321E+04-3.13634050E+01+1.58376391E+00+3.16215366E-02-1.73664942E-05    3
+4.18927663E-09-2.79899620E-13-2.12643496E+04+1.88313766E+01+0.00000000E+00    4
CH3COCH3   8/12/15      C   3H   6O   1    0G   300.000  5000.000 1394.000    21
+8.87619308E+00+1.45700263E-02-4.84823280E-06+7.38614777E-10-4.22831194E-14    2
-3.06046242E+04-2.12730484E+01+2.20008426E+00+2.74019559E-02-1.31342003E-05    3
+2.57150371E-09-6.21509091E-14-2.79933966E+04+1.55883508E+01+0.00000000E+00    4
CH3COCH2   2/14/13 THERMC   3H   5O   1    0G   300.000  5000.000 1387.000    21
+1.09524298E+01+1.11458668E-02-3.86262877E-06+6.05088857E-10-3.53293362E-14    2
-9.60833727E+03-3.15622776E+01+1.13381826E+00+3.25095045E-02-2.10424651E-05    3
+6.64421151E-09-8.12618901E-13-6.04868361E+03+2.17158655E+01+0.00000000E+00    4
CH3COCH2O2 2/14/13 THERMC   3H   5O   3    0G   300.000  5000.000 1397.000    31
+1.65756401E+01+1.06465489E-02-3.61368681E-06+5.59053564E-10-3.23832271E-14    2
-2.42541401E+04-5.45304899E+01+1.19378141E+00+4.98027161E-02-4.17999508E-05    3
+1.74527607E-08-2.88198761E-12-1.93244224E+04+2.67877493E+01+0.00000000E+00    4
CH3COCH2O  2/ 8/13 THERMC   3H   5O   2    0G   300.000  5000.000 2002.000    21
+9.84061707E+00+1.59181106E-02-5.85164644E-06+9.56160073E-10-5.75477263E-14    2
-2.11214823E+04-2.12330791E+01+5.85960137E+00+1.78954926E-02+7.41506398E-07    3
-5.40032753E-09+1.47393197E-12-1.90714739E+04+2.70987883E+00+0.00000000E+00    4
C3KET21    2/14/13 THERMC   3H   6O   3    0G   300.000  5000.000 1394.000    41
+1.75768076E+01+1.20311704E-02-4.11633942E-06+6.40149366E-10-3.72127562E-14    2
-4.15502347E+04-6.09097100E+01-8.74352903E-01+6.12501498E-02-5.51474542E-05    3
+2.48491014E-08-4.42613472E-12-3.58060819E+04+3.59306224E+01+0.00000000E+00    4
C2H3CHO           KPS12 C   3H   4O   1    0G   300.000  5000.000 1398.000    01
+9.99155394E+00+9.82348001E-03-3.31203088E-06+5.09524422E-10-2.93821890E-14    2
-1.25303509E+04-2.85168883E+01+7.33844455E-01+3.17482671E-02-2.29599468E-05    3
+8.42104232E-09-1.23613478E-12-9.38473548E+03+2.10308851E+01+0.00000000E+00    4
C2H3CO            KPS12 C   3H   3O   1    0G   300.000  5000.000 1395.000    01
+8.86032735E+00+8.48985205E-03-2.90350080E-06+4.50763986E-10-2.61524281E-14    2
+7.73489171E+03-2.06978792E+01+1.65335195E+00+2.57402596E-02-1.89009911E-05    3
+7.29174972E-09-1.16083226E-12+1.02020654E+04+1.78705872E+01+0.00000000E+00    4
C2H5CHO    8/12/15      C   3H   6O   1    0G   300.000  5000.000 1449.000    21
+1.06224453E+01+1.35569132E-02-4.60754771E-06+7.12755462E-10-4.12631683E-14    2
-2.78692266E+04-3.16628752E+01+2.18895588E+00+2.58289987E-02-6.04170058E-06    3
-3.70702654E-09+1.57131095E-12-2.42671146E+04+1.61496330E+01+0.00000000E+00    4
C2H5CO            A10/04C  3 H  5 O  1    0 G   200.000  6000.00  1000.00      1
+6.52325448E+00+1.54211952E-02-5.50898157E-06+8.85889862E-10-5.28846399E-14    2
-7.19631634E+03-5.19862218E+00+6.25722402E+00-9.17612184E-03+7.61190493E-05    3
-9.05514997E-08+3.46198215E-11-5.91616484E+03+2.23330599E+00-3.94851891E+03    4
CH2CH2CHO               C   3H   5O   1    0G   300.000  5000.000 1437.000    21
+1.00673122E+01+1.14971005E-02-3.90137798E-06+6.03029101E-10-3.48958224E-14    2
-2.75080876E+03-2.58818404E+01+2.55799036E+00+2.23391941E-02-4.89741478E-06    3
-3.58874384E-09+1.47175030E-12+4.53127696E+02+1.67016285E+01+0.00000000E+00    4
C4H10      8/12/15      C   4H  10    0    0G   300.000  5000.000 1392.000    31
+1.24923813E+01+2.15951935E-02-7.34277611E-06+1.13529859E-09-6.56730149E-14    2
-2.17598985E+04-4.41546866E+01-9.20862487E-02+4.69703816E-02-2.54761945E-05    3
+6.35894738E-09-5.16005946E-13-1.69556758E+04+2.49101571E+01+0.00000000E+00    4
PC4H9      8/12/15      C   4H   9    0    0G   300.000  5000.000 1393.000    31
+1.18547949E+01+1.96962095E-02-6.71054229E-06+1.03891144E-09-6.01513573E-14    2
+3.38182243E+03-3.72343446E+01+4.09644702E-01+4.29511341E-02-2.36582809E-05    3
+6.15744917E-09-5.64300671E-13+7.74319150E+03+2.55312526E+01+0.00000000E+00    4
SC4H9      8/12/15      C   4H   9    0    0G   300.000  5000.000 1682.000    31
+9.25139144E+00+2.24301385E-02-7.82648592E-06+1.23559460E-09-7.26249864E-14    2
+3.11148804E+03-2.16080436E+01+9.42662332E-01+3.77414530E-02-1.58911963E-05    3
+1.75489317E-09+2.89725750E-13+6.20542636E+03+2.42126605E+01+0.00000000E+00    4
PC4H9O                  C   4H   9O   1    0G   300.000  5000.000 1396.000    31
+1.53371588E+01+1.92789649E-02-6.56856538E-06+1.01724003E-09-5.89183466E-14    2
-1.41958782E+04-5.45071855E+01+1.84659093E+00+4.61054365E-02-2.44856516E-05    3
+5.11293268E-09-1.07538298E-13-9.09206746E+03+1.95237441E+01+0.00000000E+00    4
SC4H9O                  C   4H   9O   1    0G   300.000  5000.000 1411.000    31
+1.52130012E+01+1.90029969E-02-6.39004701E-06+9.80774402E-10-5.64493733E-14    2
-1.59888805E+04-5.43195369E+01+2.01772535E+00+4.70083969E-02-2.74726645E-05    3
+7.36290028E-09-6.30414237E-13-1.11892176E+04+1.74371746E+01+0.00000000E+00    4
PC4H9O2    8/12/15      C   4H   9O   2    0G   300.000  5000.000 1391.000    41
+1.66120049E+01+2.04752336E-02-7.01415262E-06+1.09010510E-09-6.32913959E-14    2
-1.57901735E+04-5.79272276E+01+1.80541406E+00+5.26493060E-02-3.30870383E-05    3
+1.04593484E-08-1.32305701E-12-1.03866773E+04+2.24829685E+01+0.00000000E+00    4
SC4H9O2                 C   4H   9O   2    0G   300.000  5000.000 1403.000    41
+1.68209433E+01+1.98834074E-02-6.71755569E-06+1.03411636E-09-5.96371075E-14    2
-1.75815350E+04-5.95731156E+01+2.27751066E+00+5.44334651E-02-3.82988187E-05    3
+1.42447767E-08-2.18864515E-12-1.25909100E+04+1.83237264E+01+0.00000000E+00    4
PC4H9O2H   8/12/15      C   4H  10O   2    0G   300.000  5000.000 1393.000    51
+1.75610913E+01+2.17832847E-02-7.46366287E-06+1.16012068E-09-6.73630029E-14    2
-3.30036118E+04-6.38547212E+01+1.04177717E+00+5.85996659E-02-3.84212378E-05    3
+1.28728231E-08-1.75491358E-12-2.70744200E+04+2.55179528E+01+0.00000000E+00    4
SC4H9O2H                C   4H  10O   2    0G   300.000  5000.000 1402.000    51
+1.78075939E+01+2.12546017E-02-7.20960281E-06+1.11291271E-09-6.43060022E-14    2
-3.48455718E+04-6.58011470E+01+1.44010868E+00+6.05300206E-02-4.36262678E-05    3
+1.66226146E-08-2.61556930E-12-2.92631492E+04+2.17354113E+01+0.00000000E+00    4
C4H8OOH1-2              C   4H   9O   2    0G   300.000  5000.000 1389.000    51
+1.67810269E+01+1.99677597E-02-6.85257220E-06+1.06628911E-09-6.19616154E-14    2
-9.14762760E+03-5.68667893E+01+2.91878364E+00+4.86143951E-02-2.81342168E-05    3
+7.64456491E-09-7.32889491E-13-3.94464787E+03+1.89326241E+01+0.00000000E+00    4
C4H8OOH1-3              C   4H   9O   2    0G   300.000  5000.000 1396.000    51
+1.61247782E+01+2.02420980E-02-6.88631475E-06+1.06534945E-09-6.16599545E-14    2
-9.16802012E+03-5.26575415E+01+2.46292502E+00+4.70131194E-02-2.42145198E-05    3
+4.65407810E-09+1.62198662E-14-3.95787917E+03+2.24569578E+01+0.00000000E+00    4
C4H8OOH1-4              C   4H   9O   2    0G   300.000  5000.000 1393.000    51
+1.69217927E+01+1.99305696E-02-6.85727522E-06+1.06879474E-09-6.21774931E-14    2
-7.87920857E+03-5.76630146E+01+1.35984095E+00+5.52812385E-02-3.75640846E-05    3
+1.32624209E-08-1.93623296E-12-2.34455867E+03+2.63197893E+01+0.00000000E+00    4
C4H8OOH2-1              C   4H   9O   2    0G   300.000  5000.000 1404.000    51
+1.77648250E+01+1.87777052E-02-6.36410476E-06+9.81958228E-10-5.67252066E-14    2
-9.93851667E+03-6.28169590E+01+2.32205003E+00+5.55032280E-02-3.97237996E-05    3
+1.47353739E-08-2.22481777E-12-4.67331585E+03+1.98332327E+01+0.00000000E+00    4
C4H8OOH2-3              C   4H   9O   2    0G   300.000  5000.000 1403.000    51
+1.70353922E+01+1.92729887E-02-6.50684653E-06+1.00126173E-09-5.77270961E-14    2
-1.09437234E+04-5.87403112E+01+3.30289851E+00+5.08231524E-02-3.39615358E-05    3
+1.17622237E-08-1.66012808E-12-6.13671017E+03+1.51726178E+01+0.00000000E+00    4
C4H8OOH2-4              C   4H   9O   2    0G   300.000  5000.000 1403.000    51
+1.72354039E+01+1.91946365E-02-6.49946502E-06+1.00210964E-09-5.78559962E-14    2
-9.71158144E+03-5.98986150E+01+1.82672511E+00+5.69912331E-02-4.24389492E-05    3
+1.67119278E-08-2.70635765E-12-4.54629884E+03+2.22051948E+01+0.00000000E+00    4
C4H8O1-2                C   4H   8O   1    0G   300.000  5000.000 1463.000    21
+1.41886108E+01+1.63162740E-02-5.16581368E-06+7.60173986E-10-4.24548403E-14    2
-2.02839382E+04-5.12817914E+01-4.29657099E+00+6.75906816E-02-5.89614134E-05    3
+2.59401158E-08-4.45926746E-12-1.48799944E+04+4.47755567E+01+0.00000000E+00    4
C4H8O1-3                C   4H   8O   1    0G   300.000  5000.000 1447.000    11
+1.32076917E+01+1.77467973E-02-5.69933762E-06+8.47771212E-10-4.77345874E-14    2
-2.11717546E+04-4.78386420E+01-5.37284363E+00+6.62224444E-02-5.35318273E-05    3
+2.19451842E-08-3.54479816E-12-1.54144887E+04+4.98345472E+01+0.00000000E+00    4
C4H8O1-4                C   4H   8O   1    0G   300.000  5000.000 1484.000    01
+1.22763349E+01+1.89105920E-02-6.09113637E-06+9.08066245E-10-5.12149503E-14    2
-2.92260872E+04-4.41235671E+01-7.78117916E+00+6.98405060E-02-5.45315920E-05    3
+2.13029617E-08-3.24666872E-12-2.28996340E+04+6.17620955E+01+0.00000000E+00    4
C4H8O2-3                C   4H   8O   1    0G   300.000  5000.000 1403.000    21
+1.06341771E+01+2.41442268E-02-1.13123977E-05+2.25480711E-09-1.54043041E-13    2
-2.10383343E+04-3.36763636E+01-4.48183187E+00+6.89313360E-02-6.15371646E-05    3
+2.73743747E-08-4.85890996E-12-1.68924193E+04+4.38882874E+01+0.00000000E+00    4
C4H8OOH1-2O2            C   4H   9O   4    0G   300.000  5000.000 1400.000    61
+2.15734750E+01+2.04528589E-02-6.99497777E-06+1.08597818E-09-6.30071127E-14    2
-2.88428166E+04-7.84560716E+01+3.02241018E+00+6.53862812E-02-4.89645658E-05    3
+1.90437784E-08-3.02309317E-12-2.25805572E+04+2.05729328E+01+0.00000000E+00    4
C4H8OOH1-3O2            C   4H   9O   4    0G   300.000  5000.000 1400.000    61
+2.15734750E+01+2.04528589E-02-6.99497777E-06+1.08597818E-09-6.30071127E-14    2
-2.88428166E+04-7.84560716E+01+3.02241018E+00+6.53862812E-02-4.89645658E-05    3
+1.90437784E-08-3.02309317E-12-2.25805572E+04+2.05729328E+01+0.00000000E+00    4
C4H8OOH1-4O2            C   4H   9O   4    0G   300.000  5000.000 1387.000    71
+2.26393370E+01+1.98017374E-02-6.92349554E-06+1.09100182E-09-6.39617643E-14    2
-2.75442161E+04-8.40747892E+01+2.91974455E+00+6.34948347E-02-4.29699499E-05    3
+1.42283155E-08-1.84506244E-12-2.04867301E+04+2.26279495E+01+0.00000000E+00    4
C4H8OOH2-1O2            C   4H   9O   4    0G   300.000  5000.000 1400.000    61
+2.15734750E+01+2.04528589E-02-6.99497777E-06+1.08597818E-09-6.30071127E-14    2
-2.88428166E+04-7.84560716E+01+3.02241018E+00+6.53862812E-02-4.89645658E-05    3
+1.90437784E-08-3.02309317E-12-2.25805572E+04+2.05729328E+01+0.00000000E+00    4
C4H8OOH2-3O2            C   4H   9O   4    0G   300.000  5000.000 1408.000    61
+2.19463055E+01+1.97307584E-02-6.65765380E-06+1.02424556E-09-5.90486257E-14    2
-3.07772334E+04-8.12053531E+01+3.34683971E+00+6.67468082E-02-5.25088611E-05    3
+2.14288389E-08-3.53381793E-12-2.47340662E+04+1.73189003E+01+0.00000000E+00    4
C4H8OOH2-4O2            C   4H   9O   4    0G   300.000  5000.000 1400.000    61
+2.15734750E+01+2.04528589E-02-6.99497777E-06+1.08597818E-09-6.30071127E-14    2
-2.88428166E+04-7.84560716E+01+3.02241018E+00+6.53862812E-02-4.89645658E-05    3
+1.90437784E-08-3.02309317E-12-2.25805572E+04+2.05729328E+01+0.00000000E+00    4
C4H71-2,4OOH            C   4H   9O   4    0G   300.000  5000.000 1398.000    71
+2.18629952E+01+1.99359398E-02-6.85103949E-06+1.06712096E-09-6.20561893E-14    2
-2.10042547E+04-7.80706874E+01+2.99387028E+00+6.52913914E-02-4.87958562E-05    3
+1.88107554E-08-2.95256716E-12-1.46021097E+04+2.27763716E+01+0.00000000E+00    4
C4H72-1,3OOH            C   4H   9O   4    0G   300.000  5000.000 1395.000    71
+2.14626449E+01+2.02946207E-02-6.97889021E-06+1.08750673E-09-6.32605387E-14    2
-2.22196721E+04-7.60671568E+01+3.85542428E+00+6.05523559E-02-4.18122063E-05    3
+1.46680029E-08-2.07881996E-12-1.60359412E+04+1.87734959E+01+0.00000000E+00    4
C4H72-1,4OOH            C   4H   9O   4    0G   300.000  5000.000 1387.000    71
+2.10228668E+01+2.10127561E-02-7.30349553E-06+1.14623341E-09-6.70076491E-14    2
-2.02908167E+04-7.29927491E+01+3.41714555E+00+5.89885977E-02-3.76843121E-05    3
+1.18450422E-08-1.46347291E-12-1.38437952E+04+2.27094787E+01+0.00000000E+00    4
C4H71-2,3OOH            C   4H   9O   4    0G   300.000  5000.000 1406.000    71
+2.22828679E+01+1.92253507E-02-6.52860872E-06+1.00881573E-09-5.83408336E-14    2
-2.29719991E+04-8.11231836E+01+3.30790561E+00+6.66513240E-02-5.21744859E-05    3
+2.10434152E-08-3.42495389E-12-1.67536738E+04+1.95806784E+01+0.00000000E+00    4
C4H7O1-3OOH-4           C   4H   8O   3    0G   300.000  5000.000 1418.000    31
+1.87250111E+01+1.88463312E-02-6.40165949E-06+9.89754621E-10-5.72727585E-14    2
-3.29825730E+04-7.18225468E+01-5.40949665E+00+8.05102667E-02-6.64646030E-05    3
+2.73711905E-08-4.44856733E-12-2.53005240E+04+5.56327196E+01+0.00000000E+00    4
C4H7O1-3OOH-2           C   4H   8O   3    0G   300.000  5000.000 1425.000    31
+1.97110479E+01+1.79060432E-02-6.05724664E-06+9.34110479E-10-5.39628469E-14    2
-3.52532541E+04-7.83129016E+01-4.68244067E+00+8.03419743E-02-6.67264700E-05    3
+2.74081300E-08-4.41623778E-12-2.75307409E+04+5.04193128E+01+0.00000000E+00    4
C4H7O1-2OOH-4           C   4H   8O   3    0G   300.000  5000.000 1417.000    41
+1.96187267E+01+1.77382423E-02-6.03563743E-06+9.34268374E-10-5.41073277E-14    2
-3.21917914E+04-7.50295988E+01-3.06056578E+00+7.52777235E-02-6.16382083E-05    3
+2.51520765E-08-4.05109146E-12-2.49310387E+04+4.48871201E+01+0.00000000E+00    4
C4H7O1-4OOH-2           C   4H   8O   3    0G   300.000  5000.000 1470.000    21
+1.74906412E+01+1.87794733E-02-6.05491558E-06+9.03185679E-10-5.09571870E-14    2
-4.22716632E+04-6.51860330E+01-5.17426936E+00+7.89225917E-02-6.62654132E-05    3
+2.77698767E-08-4.54377840E-12-3.53780833E+04+5.35508489E+01+0.00000000E+00    4
C4H7O1-2OOH-3           C   4H   8O   3    0G   300.000  5000.000 1435.000    41
+1.83476383E+01+1.72627711E-02-5.53440131E-06+8.21396496E-10-4.61479654E-14    2
-3.29223599E+04-6.69919656E+01-9.44964311E-01+7.31026695E-02-6.71227799E-05    3
+3.12252290E-08-5.67206759E-12-2.74510619E+04+3.25427282E+01+0.00000000E+00    4
C4H7O2-3OOH-1           C   4H   8O   3    0G   300.000  5000.000 1424.000    41
+2.03028185E+01+1.69331534E-02-5.71128715E-06+8.79005552E-10-5.07088176E-14    2
-3.43451470E+04-7.95919117E+01-3.04171082E+00+7.75254740E-02-6.55776743E-05    3
+2.74944445E-08-4.52476822E-12-2.70343494E+04+4.33136810E+01+0.00000000E+00    4
C4H72-1OOH              C   4H   8O   2    0G   300.000  5000.000 1381.000    41
+1.80122740E+01+1.70340943E-02-5.89884086E-06+9.23962123E-10-5.39539803E-14    2
-1.74585465E+04-6.55209757E+01+1.29755275E+00+5.59252255E-02-4.08890003E-05    3
+1.54880526E-08-2.42412478E-12-1.16046928E+04+2.43621382E+01+0.00000000E+00    4
NC4KET12                C   4H   8O   3    0G   300.000  5000.000 1389.000    51
+2.17577434E+01+1.64473301E-02-5.79961988E-06+9.19149624E-10-5.41037382E-14    2
-4.47115295E+04-8.37725285E+01-7.24231793E-01+7.26648886E-02-6.04779190E-05    3
+2.54348857E-08-4.30152907E-12-3.72936909E+04+3.56276963E+01+0.00000000E+00    4
NC4KET13                C   4H   8O   3    0G   300.000  5000.000 1411.000    51
+1.93085398E+01+1.73455091E-02-5.85046818E-06+9.00297947E-10-5.19274609E-14    2
-4.51023813E+04-7.04869509E+01+3.31775682E+00+5.28482064E-02-3.43211665E-05    3
+1.04562704E-08-1.12796519E-12-3.94868388E+04+1.58443308E+01+0.00000000E+00    4
NC4KET14                C   4H   8O   3    0G   300.000  5000.000 1385.000    51
+1.89231898E+01+1.82270124E-02-6.27434124E-06+9.78729382E-10-5.69844333E-14    2
-4.32508875E+04-6.78717188E+01+2.92378737E+00+5.07578011E-02-2.88360718E-05    3
+6.64649914E-09-2.83907499E-13-3.72946444E+04+1.96328202E+01+0.00000000E+00    4
NC4KET21                C   4H   8O   3    0G   300.000  5000.000 1389.000    51
+2.10786402E+01+1.61788162E-02-5.53076294E-06+8.59641186E-10-4.99535144E-14    2
-4.57563821E+04-7.88014765E+01-3.88449068E-01+6.92735051E-02-5.58731127E-05    3
+2.25791086E-08-3.63900158E-12-3.86875801E+04+3.52948090E+01+0.00000000E+00    4
NC4KET23                C   4H   8O   3    0G   300.000  5000.000 1411.000    51
+1.76877593E+01+1.84820224E-02-6.18384585E-06+9.45792334E-10-5.42981801E-14    2
-4.78594254E+04-6.06681612E+01+3.56926969E+00+5.20285891E-02-3.64134216E-05    3
+1.32007682E-08-1.93576774E-12-4.30650503E+04+1.48669401E+01+0.00000000E+00    4
NC4KET24                C   4H   8O   3    0G   300.000  5000.000 1394.000    51
+1.74146206E+01+1.92744267E-02-6.57971403E-06+1.02023879E-09-5.91418353E-14    2
-4.60663138E+04-5.80320911E+01+3.12062686E+00+5.01343936E-02-3.10194950E-05    3
+9.36512355E-09-1.07548923E-12-4.08644270E+04+1.96071994E+01+0.00000000E+00    4
C4H71-3OOH              C   4H   8O   2    0G   300.000  5000.000 1392.000    41
+1.92985494E+01+1.54534427E-02-5.25460431E-06+8.13772446E-10-4.71689947E-14    2
-1.85003480E+04-7.49926639E+01-1.50977396E+00+6.85369305E-02-5.75193633E-05    3
+2.43179107E-08-4.09788488E-12-1.18018961E+04+3.50420113E+01+0.00000000E+00    4
C4H71-4OOH              C   4H   8O   2    0G   300.000  5000.000 1392.000    41
+1.59871304E+01+1.86028119E-02-6.40003189E-06+9.97531711E-10-5.80334203E-14    2
-1.70152141E+04-5.46227137E+01+1.31653247E+00+5.16546159E-02-3.47310922E-05    3
+1.20405755E-08-1.71650639E-12-1.17754576E+04+2.46384545E+01+0.00000000E+00    4
C4H71-3,4OOH            C   4H   9O   4    0G   300.000  5000.000 1400.000    71
+2.18394783E+01+1.98802807E-02-6.81505369E-06+1.05975117E-09-6.15560073E-14    2
-2.09468667E+04-7.79984909E+01+2.56890026E+00+6.71962184E-02-5.16999792E-05    3
+2.05770379E-08-3.32914310E-12-1.45125600E+04+2.46332539E+01+0.00000000E+00    4
C4H72-3,4OOH            C   4H   9O   4    0G   300.000  5000.000 1395.000    71
+2.14626449E+01+2.02946207E-02-6.97889021E-06+1.08750673E-09-6.32605387E-14    2
-2.22196721E+04-7.60671568E+01+3.85542428E+00+6.05523559E-02-4.18122063E-05    3
+1.46680029E-08-2.07881996E-12-1.60359412E+04+1.87734959E+01+0.00000000E+00    4
HO2CH2CHO  9/ 8/14      C   2H   4O   3    0G   300.000  5000.000 1391.000    31
+1.51554685E+01+7.57240000E-03-2.72693024E-06+4.38217189E-10-2.60434287E-14    2
-3.41419680E+04-5.01255068E+01-1.32768631E+00+5.21618601E-02-4.97327645E-05    3
+2.31272366E-08-4.20787867E-12-2.90608844E+04+3.61860491E+01+0.00000000E+00    4
C4H71-O   11/13/18 THERMC   4H   7O   1    0G   300.000  5000.000 1369.000    21 !UB REFIT 13-11-2018
 1.56996664E+01 1.61014619E-02-6.49436831E-06 1.11548710E-09-6.91568286E-14    2
-1.62497835E+03-5.78467858E+01 6.10872657E+00 2.28749673E-02 3.92794486E-06    3
-1.04315787E-08 2.89510888E-12 3.53302055E+03-3.49511801E-01                   4
IC4H10     8/12/15      C   4H  10    0    0G   300.000  5000.000 1397.000    31
+1.26422737E+01+2.14133551E-02-7.26711536E-06+1.12207226E-09-6.48434177E-14    2
-2.28293782E+04-4.66059659E+01-1.07413829E+00+5.24618320E-02-3.42407949E-05    3
+1.18817533E-08-1.73238254E-12-1.79218932E+04+2.74851665E+01+0.00000000E+00    4
IC4H9      8/12/15      C   4H   9    0    0G   300.000  5000.000 1397.000    31
+1.23261837E+01+1.92057770E-02-6.52063623E-06+1.00704497E-09-5.82038734E-14    2
+2.50995714E+03-4.13478742E+01+1.20802408E-01+4.73187324E-02-3.16440251E-05    3
+1.14229699E-08-1.74784642E-12+6.84032915E+03+2.44291032E+01+0.00000000E+00    4
TC4H9      8/12/15      C   4H   9    0    0G   300.000  5000.000 1380.000    31
+1.02682832E+01+2.09965262E-02-7.14945754E-06+1.10648358E-09-6.40498314E-14    2
+1.57542675E+02-3.00960941E+01+1.05841769E+00+3.41133739E-02-9.03156779E-06    3
-2.95313136E-09+1.41436845E-12+4.22699258E+03+2.23965051E+01+0.00000000E+00    4
TC4H9O            T08/04C  4 H  9 O  1    0 G   200.000  6000.00  1000.00      1
+1.27371509E+01+2.33707342E-02-8.50516678E-06+1.38519973E-09-8.34398061E-14    2
-1.66940150E+04-4.53156321E+01+2.77057100E+00+2.68033175E-02+4.12718360E-05    3
-7.22054739E-08+3.02642276E-11-1.27079262E+04+1.21532856E+01-1.04543262E+04    4
IC4H9O            A08/04C  4 H  9 O  1    0 G   200.000  6000.00  1000.00      1
+1.16309708E+01+2.47981574E-02-9.01550536E-06+1.46714720E-09-8.83214518E-14    2
-1.37854612E+04-3.81956151E+01+3.80297372E+00+1.56874209E-02+6.81105412E-05    3
-9.83346774E-08+3.95261902E-11-1.00832243E+04+9.78963305E+00-7.82602559E+03    4
IC3H7CHO   2/22/96 THERMC   4H   8O   1    0G   300.000  5000.000 1391.000    31
+1.37501656E+01+1.83126722E-02-6.28572629E-06+9.78250756E-10-5.68538653E-14    2
-3.26936771E+04-4.77270548E+01-2.73021382E-01+4.89696307E-02-3.12770049E-05    3
+1.00052945E-08-1.27512074E-12-2.76054737E+04+2.83451139E+01+0.00000000E+00    4
SC4H7OH-I         L 2/00C   4H   8O   1    0G   300.000  5000.000 1395.000    31
+1.30299481E+01+1.83782479E-02-6.18529878E-06+9.49578099E-10-5.46526348E-14    2
-3.10723026E+04-4.22891828E+01+2.70103499E+00+4.17950180E-02-2.67860575E-05    3
+9.38191037E-09-1.41171285E-12-2.73561190E+04+1.35316306E+01+0.00000000E+00    4
IC4H6OH                 C   4H   7O   1    0G   300.000  5000.000 1402.000    21
+1.53490714E+01+1.38856699E-02-4.56427754E-06+6.90418690E-10-3.93540403E-14    2
-1.20164758E+04-5.55975530E+01-1.46664187E+00+6.03351671E-02-5.43112644E-05    3
+2.49299933E-08-4.52282491E-12-6.95012413E+03+3.20768458E+01+0.00000000E+00    4
IC3H7CO    2/22/96 THERMC   4H   7O   1    0G   300.000  5000.000 1390.000    31
+1.33305736E+01+1.61873930E-02-5.56711402E-06+8.67575951E-10-5.04696549E-14    2
-1.37307001E+04-4.33958746E+01+5.03452639E-01+4.41607510E-02-2.82139091E-05    3
+8.93548675E-09-1.11327422E-12-9.07755468E+03+2.61991461E+01+0.00000000E+00    4
IC3H6CHO   2/22/96 THERMC   4H   7O   1    0G   300.000  5000.000 1390.000    31
+1.33102250E+01+1.62097959E-02-5.57575891E-06+8.69003718E-10-5.05554202E-14    2
-7.62177931E+03-4.25050854E+01+5.21481767E-01+4.43114357E-02-2.86617314E-05    3
+9.30319894E-09-1.20761563E-12-2.99677086E+03+2.68182130E+01+0.00000000E+00    4
TC3H6CHO   2/22/96 THERMC   4H   7O   1    0G   300.000  5000.000 1389.000    21
+1.31013047E+01+1.66391865E-02-5.68457623E-06+8.81808351E-10-5.11290161E-14    2
-1.30638647E+04-4.42705813E+01+1.87052762E+00+4.14869677E-02-2.66815701E-05    3
+9.01531610E-09-1.27870633E-12-8.97730744E+03+1.66174178E+01+0.00000000E+00    4
IC3H5CHO                C   4H   6O   1    0G   300.000  5000.000 1396.000    21
+1.33892118E+01+1.39115420E-02-4.75820958E-06+7.38736618E-10-4.28606559E-14    2
-1.97917448E+04-4.60146004E+01+1.09372823E+00+4.43315368E-02-3.41918451E-05    3
+1.39369607E-08-2.33791460E-12-1.56745978E+04+1.94458467E+01+0.00000000E+00    4
IC3H6CO   03/03/95 THERMC   4H   6O   1    0G   300.000  5000.000 1397.00     41
+1.32548232E+01+1.40142787E-02-4.78910215E-06+7.42924342E-10-4.30737566E-14    2
-2.00529779E+04-4.44810221E+01+2.28039055E+00+4.17016989E-02-3.25089661E-05    3
+1.37243419E-08-2.40573132E-12-1.63939712E+04+1.38187714E+01+0.00000000E+00    4
IC3H5CO                 C   4H   5O   1    0G   300.000  5000.000 1396.000    21
+1.29634401E+01+1.17954996E-02-4.04361488E-06+6.28771516E-10-3.65209867E-14    2
-8.26519462E+02-4.20562575E+01+1.87306990E+00+3.95188508E-02-3.11404053E-05    3
+1.28844447E-08-2.18165308E-12+2.85270691E+03+1.68774016E+01+0.00000000E+00    4
IC3H4CHO-A              C   4H   5O   1    0G   300.000  5000.000 1392.000    11
+1.41736959E+01+1.09161978E-02-3.69020878E-06+5.69228087E-10-3.29023246E-14    2
-1.92867979E+03-5.02663740E+01+7.64345054E-01+4.45242412E-02-3.61033720E-05    3
+1.48295287E-08-2.43809290E-12+2.44732544E+03+2.08541848E+01+0.00000000E+00    4
IC4H8O     9/ 1/12      C   4H   8O   1    0G   300.000  5000.000 1394.000    21
+1.40433578E+01+2.05733637E-02-9.09519220E-06+1.73417298E-09-1.14908544E-13    2
-3.62275308E+04-6.90009668E+01-5.02573822E+00+7.51340960E-02-6.88668822E-05    3
+3.12223247E-08-5.60128818E-12-3.07481413E+04+2.96284295E+01+0.00000000E+00    4
TC3H6O2CHO 8/ 2/95 THERMC   4H   7O   3    0G   300.000  5000.000 1386.00     41
+1.85534443E+01+1.68774389E-02-5.90752965E-06+9.31518085E-10-5.46345187E-14    2
-2.85447191E+04-6.82486667E+01+2.17883383E+00+5.41595832E-02-3.83435886E-05    3
+1.38308104E-08-2.04190147E-12-2.27394154E+04+2.00751264E+01+0.00000000E+00    4
IC3H5O2HCHO 8/2/95 THERMC   4H   7O   3    0G   300.000  5000.000 1387.00     51
+2.06288832E+01+1.48625539E-02-5.25305276E-06+8.33772951E-10-4.91277401E-14    2
-2.27589076E+04-7.82962888E+01+2.05984770E+00+5.82331716E-02-4.37672100E-05    3
+1.63249918E-08-2.43462051E-12-1.63496250E+04+2.13687921E+01+0.00000000E+00    4
TC3H6O2HCO 8/ 2/95 THERMC   4H   7O   3    0G   300.000  5000.000 1387.00     51
+2.06472678E+01+1.48526500E-02-5.25104875E-06+8.33619219E-10-4.91256069E-14    2
-2.88719869E+04-7.95951389E+01+2.03864428E+00+5.80421003E-02-4.32123528E-05    3
+1.58792094E-08-2.32209543E-12-2.24284673E+04+2.03680990E+01+0.00000000E+00    4
TC3H6OCHO  8/25/95 THERMC   4H   7O   2    0G   300.000  5000.000 1394.00     31
+1.70371287E+01+1.54400645E-02-5.28332886E-06+8.21085347E-10-4.76898429E-14    2
-2.75871941E+04-6.37271230E+01+3.70830259E-01+5.38475661E-02-3.82477565E-05    3
+1.32882237E-08-1.79228730E-12-2.18391262E+04+2.58142112E+01+0.00000000E+00    4
IC4H9O2    9/ 1/12      C   4H   9O   2    0G   300.000  5000.000 1432.000    41
+1.78793870E+01+1.82474607E-02-6.01252193E-06+9.11106794E-10-5.20018932E-14    2
-1.74569774E+04-6.61552973E+01+1.77219624E+00+5.34032789E-02-3.31041810E-05    3
+9.24465657E-09-8.01706642E-13-1.17768774E+04+2.09581481E+01+0.00000000E+00    4
TC4H9O2    9/ 1/12      C   4H   9O   2    0G   300.000  5000.000 1380.000    41
+1.80863238E+01+1.99282971E-02-6.98287309E-06+1.10171726E-09-6.46381057E-14    2
-2.04420664E+04-6.97533212E+01+2.63892371E+00+5.44717499E-02-3.75504698E-05    3
+1.40479250E-08-2.27968600E-12-1.47598933E+04+1.40325533E+01+0.00000000E+00    4
IC4H8O2H-I 9/ 1/12      C   4H   9O   2    0G   300.000  5000.000 1414.000    51
+1.83915486E+01+1.73042831E-02-5.66841018E-06+8.55414265E-10-4.86781778E-14    2
-9.48569748E+03-6.67673286E+01+1.86432620E-01+6.26430177E-02-4.83690886E-05    3
+1.88657148E-08-2.91189385E-12-3.59086611E+03+2.97635367E+01+0.00000000E+00    4
IC4H8O2H-T 9/ 1/12      C   4H   9O   2    0G   300.000  5000.000 1413.000    51
+1.69753885E+01+1.85198010E-02-6.09075415E-06+9.21673609E-10-5.25502501E-14    2
-1.14812757E+04-5.88259039E+01+3.84374544E+00+4.36800978E-02-2.07599526E-05    3
+2.51709167E-09+5.41306513E-13-6.50766215E+03+1.34244877E+01+0.00000000E+00    4
TC4H8O2H-I 9/ 1/12      C   4H   9O   2    0G   300.000  5000.000 1379.000    51
+1.81415374E+01+1.94699499E-02-6.82750014E-06+1.07773311E-09-6.32519099E-14    2
-1.23570939E+04-6.63491602E+01+3.54378349E+00+5.25201369E-02-3.69898493E-05    3
+1.44634925E-08-2.47536050E-12-6.98183185E+03+1.27623539E+01+0.00000000E+00    4
CC4H8O     9/ 1/12      C   4H   8O   1    0G   300.000  5000.000 1431.000    11
+1.51841776E+01+1.64656666E-02-5.33483091E-06+7.98149768E-10-4.51160381E-14    2
-3.33923434E+04-7.43746988E+01-6.56746688E+00+7.87298554E-02-7.33065478E-05    3
+3.40602701E-08-6.15674656E-12-2.71582518E+04+3.80875851E+01+0.00000000E+00    4
IC4H8OOH-IO2 9/ 1/12    C   4H   9O   4    0G   300.000  5000.000 1367.000    61
+2.24664901E+01+2.09351287E-02-7.44324128E-06+1.18589255E-09-7.00546897E-14    2
-2.94495457E+04-8.54241451E+01+4.23354857E+00+5.63088857E-02-3.15672522E-05    3
+7.79536931E-09-6.21665008E-13-2.22782534E+04+1.52623111E+01+0.00000000E+00    4
IC4H8OOH-TO2 9/ 1/12    C   4H   9O   4    0G   300.000  5000.000 1385.000    61
+2.32464612E+01+1.88384513E-02-6.40938087E-06+9.92649459E-10-5.75275879E-14    2
-3.16533132E+04-8.88301710E+01+3.36413530E+00+6.93742776E-02-5.70416393E-05    3
+2.46040165E-08-4.32848680E-12-2.51137558E+04+1.65767339E+01+0.00000000E+00    4
TC4H8OOH-IO2 9/ 1/12    C   4H   9O   4    0G   300.000  5000.000 1385.000    61
+2.32464612E+01+1.88384513E-02-6.40938087E-06+9.92649459E-10-5.75275879E-14    2
-3.16533132E+04-8.88301710E+01+3.36413530E+00+6.93742776E-02-5.70416393E-05    3
+2.46040165E-08-4.32848680E-12-2.51137558E+04+1.65767339E+01+0.00000000E+00    4
IC4KETII   7/19/ 0 THERMC   4H   8O   3    0G   300.000  5000.000 1387.000    51
+1.95143059E+01+1.82377395E-02-6.38908606E-06+1.00801571E-09-5.91440350E-14    2
-4.46884836E+04-7.17167584E+01+1.15501614E+00+6.10622345E-02-4.49711323E-05    3
+1.70514654E-08-2.65948602E-12-3.82747956E+04+2.69612235E+01+0.00000000E+00    4
IC4KETIT   7/19/ 0 THERMC   4H   8O   3    0G   300.000  5000.000 1388.000    51
+2.09369850E+01+1.71090955E-02-6.01892169E-06+9.52353863E-10-5.59926176E-14    2
-4.77819819E+04-8.27717611E+01+1.14243741E+00+6.33840797E-02-4.73084738E-05    3
+1.77145373E-08-2.67265475E-12-4.09366796E+04+2.34844867E+01+0.00000000E+00    4
TIC4H7Q2-I 5/ 6/96 THERMC   4H   9O   4    0G   300.000  5000.000 1400.000    71
+2.33848631E+01+1.87070035E-02-6.44021945E-06+1.00428123E-09-5.84468189E-14    2
-2.61180902E+04-8.76610135E+01+4.48426361E+00+6.61225007E-02-5.27349018E-05    3
+2.18215585E-08-3.66788946E-12-1.98906586E+04+1.26719614E+01+0.00000000E+00    4
IIC4H7Q2-I 7/15/96 THERMC   4H   9O   4    0G   300.000  5000.000 1394.000    71
+2.30500244E+01+1.92149194E-02-6.66622576E-06+1.04495725E-09-6.10370520E-14    2
-2.32086881E+04-8.39949885E+01+4.93055661E+00+6.05819201E-02-4.23665566E-05    3
+1.49122008E-08-2.10978665E-12-1.68415495E+04+1.36228018E+01+0.00000000E+00    4
IIC4H7Q2-T 7/15/96 THERMC   4H   9O   4    0G   300.000  5000.000 1377.000    71
+2.15070321E+01+2.05359839E-02-7.12383399E-06+1.11655053E-09-6.52112103E-14    2
-2.51117508E+04-7.43379783E+01+8.16274487E+00+4.34463050E-02-1.76972456E-05    3
+4.88790666E-10+9.03915465E-13-1.96501749E+04+2.62067299E-01+0.00000000E+00    4
IC4H7OOH   4/15/15      C   4H   8O   2    0G   300.000  5000.000 1386.000    41
+1.82897194E+01+1.67815784E-02-5.80668193E-06+9.08949180E-10-5.30513302E-14    2
-1.82046522E+04-6.72111342E+01+1.31851762E-01+6.19561224E-02-4.99343877E-05    3
+2.09628211E-08-3.59717924E-12-1.21399925E+04+2.93905962E+01+0.00000000E+00    4
IC4H9O2H   9/ 1/12      C   4H  10O   2    0G   300.000  5000.000 1402.000    51
+1.91651624E+01+1.93678648E-02-6.41984435E-06+9.76947752E-10-5.59299558E-14    2
-3.48790978E+04-7.42063787E+01-5.47969191E-01+6.57428787E-02-4.70123149E-05    3
+1.65991096E-08-2.27331437E-12-2.82180462E+04+3.12961385E+01+0.00000000E+00    4
TC4H9O2H   9/ 1/12      C   4H  10O   2    0G   300.000  5000.000 1382.000    51
+1.90926853E+01+2.12697804E-02-7.46252626E-06+1.17841127E-09-6.91795087E-14    2
-3.77278405E+04-7.61321196E+01+4.45573540E-01+6.66153523E-02-5.20932123E-05    3
+2.22301799E-08-4.00189859E-12-3.12260714E+04+2.37278262E+01+0.00000000E+00    4
IC4H8      8/12/15      C   4H   8    0    0G   300.000  5000.000 1392.000    21
+1.11444028E+01+1.81609265E-02-6.17791116E-06+9.55481871E-10-5.52826092E-14    2
-7.84024684E+03-3.68508829E+01+5.72478139E-02+4.17768938E-02-2.49095729E-05    3
+7.54294402E-09-9.23202212E-13-3.72166259E+03+2.35698905E+01+0.00000000E+00    4
IC4H7      8/12/15      C   4H   7    0    0G   300.000  5000.000 1384.000    11
+1.18999143E+01+1.51569859E-02-5.09995449E-06+7.83722199E-10-4.51660275E-14    2
+1.00363555E+04-4.02286635E+01-2.29578762E-01+4.17842986E-02-2.66885700E-05    3
+8.42205744E-09-1.03175361E-12+1.43946680E+04+2.54797645E+01+0.00000000E+00    4
IC4H7-I1   5/13/15      C   4H   7    0    0G   300.000  5000.000 1396.000    21
+1.11158752E+01+1.55127192E-02-5.23769366E-06+8.05998394E-10-4.64703390E-14    2
+2.19488297E+04-3.41440480E+01+9.12464579E-01+3.88654394E-02-2.57575714E-05    3
+9.07760026E-09-1.33946902E-12+2.55635553E+04+2.08634918E+01+0.00000000E+00    4
IC4H7O2           L 2/00C   4H   7O   2    0G   300.000  5000.000 1404.000    31
+1.45791608E+01+1.62136068E-02-5.26957103E-06+7.90454323E-10-4.47755051E-14    2
-1.20848042E+03-4.56459433E+01+1.43532045E+00+4.89026570E-02-3.63600970E-05    3
+1.41906420E-08-2.24557878E-12+3.09284623E+03+2.41320196E+01+0.00000000E+00    4
IC4H6OOH-I        L 2/00C   4H   7O   2    0G   300.000  5000.000 1398.000    31
+1.73601429E+01+1.42046196E-02-4.65348263E-06+7.02209785E-10-3.99552775E-14    2
-1.07509366E+03-6.12822377E+01+6.06669321E+00+3.94950065E-02-2.52721718E-05    3
+7.84485641E-09-8.98876886E-13+2.87448422E+03-3.78377026E-01+0.00000000E+00    4
CCYCCOOC-T1        THERMC   4H   7O   2    0G   300.000  5000.000 1394.000    11
+1.68269657E+01+1.64471921E-02-5.63767184E-06+8.78001611E-10-5.10959632E-14    2
-3.65710841E+03-6.74096786E+01-5.29767923E+00+6.65082201E-02-4.67054235E-05    3
+1.51029775E-08-1.74322091E-12+3.97935712E+03+5.16412476E+01+0.00000000E+00    4
C2CYCOOC-I1   7/14      C   4H   7O   2    0G   300.000  5000.000 1388.000    21
+1.89745085E+01+1.50113808E-02-5.30728309E-06+8.42454740E-10-4.96392976E-14    2
-6.93111358E+03-9.08581019E+01-2.04718031E+00+7.26608379E-02-6.82960279E-05    3
+3.27505762E-08-6.23802161E-12-3.71475599E+02+1.92056057E+01+0.00000000E+00    4
CCYCCOOC-I2       L 2/00C   4H   7O   2    0G   300.000  5000.000 1398.000    11
+1.63388791E+01+1.65879474E-02-5.61829108E-06+8.67331033E-10-5.01476782E-14    2
+6.66946988E+03-6.40322040E+01-4.55772603E+00+7.10221387E-02-6.05228430E-05    3
+2.61773944E-08-4.51390528E-12+1.32922215E+04+4.60828737E+01+0.00000000E+00    4
IC3H5OOCH2        L 2/00C   4H   7O   2    0G   300.000  5000.000 1410.000    41
+5.05335676E+00+3.62904388E-02-1.54012992E-05+2.74341619E-09-1.74718602E-13    2
+4.08326144E+03-2.55389509E+00-1.26548168E+00-3.61337863E-03+7.31803998E-05    3
-5.49845697E-08+1.20447492E-11+1.33108969E+04+5.33428723E+01+0.00000000E+00    4
CHOIC3H6O         L 2/00C   4H   7O   2    0G   300.000  5000.000 1386.000    31
+1.55511970E+01+1.67360034E-02-5.73573457E-06+8.92095191E-10-5.18351848E-14    2
-2.50674335E+04-5.23215658E+01+2.55559437E-01+5.22086026E-02-3.72283766E-05    3
+1.36714420E-08-2.05638885E-12-1.97284649E+04+2.99210251E+01+0.00000000E+00    4
CVCYCCOC          L 2/00C   4H   6O   1    0G   300.000  5000.000 1397.000     1
+1.14363523E+01+1.63250968E-02-5.57146218E-06+8.63795613E-10-5.00701899E-14    2
-5.44653450E+03-3.87179379E+01-2.45566808E+00+4.88377067E-02-3.46186324E-05    3
+1.26590643E-08-1.88737988E-12-6.43460880E+02+3.58434061E+01+0.00000000E+00    4
CCYC2OCO          L 2/00C   4H   7O   2    0G   300.000  5000.000 1401.000    21
+1.64352871E+01+1.65843210E-02-5.71790511E-06+8.92586562E-10-5.19865043E-14    2
-1.60938498E+04-5.96946106E+01-2.97381263E+00+6.75615160E-02-5.79901709E-05    3
+2.55213006E-08-4.49991674E-12-9.93607156E+03+4.25127997E+01+0.00000000E+00    4
CCYCCO-T1         L 2/00C   3H   5O   1    0G   300.000  5000.000 1389.000    11
+1.03394781E+01+1.15180335E-02-3.87496644E-06+5.95744364E-10-3.43539552E-14    2
+7.17658970E+03-2.89687593E+01-1.39311392E+00+3.81789194E-02-2.62316288E-05    3
+8.74877238E-09-1.11296763E-12+1.12534953E+04+3.41877003E+01+0.00000000E+00    4
IC4H7O     4/ 3/ 0 THERMC   4H   7O   1    0G   300.000  5000.000 1386.000    21
+1.33457615E+01+1.61218588E-02-5.44376403E-06+8.38199374E-10-4.83608280E-14    2
+6.11443644E+02-4.36818838E+01+1.74700687E+00+4.07783436E-02-2.44750243E-05    3
+7.06502958E-09-7.51570589E-13+4.86979233E+03+1.94535999E+01+0.00000000E+00    4
IC3H5OCH2  6/ 2/14 CZHOUH   7C   4O   1     G   298.150  2000.000 1000.00      1
+6.64731727E+00+3.08190709E-02-1.73209320E-05+5.01099629E-09-6.00089387E-13    2
+1.70679921E+03-5.91214819E+00-2.14798958E+00+7.00225553E-02-8.21595440E-05    3
+5.22589946E-08-1.34176532E-11+3.26474773E+03+3.55145589E+01+0.00000000E+00    4
IC4H7OOCH3              C   5H  10O   2    0G   300.000  5000.000 1386.000    51
+1.95896715E+01+2.31057369E-02-8.02911330E-06+1.25969946E-09-7.36169360E-14    2
-1.80069088E+04-7.34192482E+01+1.26784161E+00+6.82442475E-02-5.30807931E-05    3
+2.27496198E-08-4.11475065E-12-1.16767937E+04+2.44900544E+01+0.00000000E+00    4
IC4H7OOIC4H7            C   8H  14O   2    0G   300.000  5000.000 1390.000    71
+2.80447245E+01+3.27505220E-02-1.13220177E-05+1.77027767E-09-1.03211988E-13    2
-1.72683337E+04-1.15134796E+02-2.07881710E-01+1.04075647E-01-8.33973077E-05    3
+3.60897624E-08-6.47906520E-12-7.79062693E+03+3.50446555E+01+0.00000000E+00    4
C4H8-1                  C   4H   8    0    0G   300.000  5000.000 1388.000    21
+1.10189295E+01+1.82714177E-02-6.21801907E-06+9.62038611E-10-5.56791341E-14    2
-5.80998818E+03-3.47942287E+01+1.62599556E-01+4.01052746E-02-2.18038592E-05    3
+5.47070727E-09-4.54073315E-13-1.65402601E+03+2.48169258E+01+0.00000000E+00    4
C4H71-1                 H   7C   4          G   298.150  2000.000 1000.00      1 !CWZ ADDED FROM YL CALCULATION
+4.93165379E+00+2.62974295E-02-1.16478367E-05+2.24008697E-09-1.22866440E-13    2
+2.68061697E+04+1.40495737E+00+1.73186779E+00+3.50026587E-02-1.85648084E-05    3
+2.75748675E-09+7.71262301E-13+2.76508226E+04+1.78655539E+01+0.00000000E+00    4
C4H71-1                 C   4H   7    0    0G   300.000  5000.000 1390.000    21
+1.10531750E+01+1.55668782E-02-5.25853044E-06+8.09627095E-10-4.67015477E-14    2
+2.39455759E+04-3.31548457E+01+8.97231085E-01+3.77003788E-02-2.33194855E-05    3
+7.38468124E-09-9.50027900E-13+2.76498158E+04+2.19835413E+01+0.00000000E+00    4
C4H71-2                 H   7C   4          G   298.150  2000.000 1000.00      1 !CWZ ADDED FROM YL CALCULATION
+4.57642739E+00+2.64291321E-02-1.13345708E-05+1.98119158E-09-6.72515039E-14    2
+2.51643094E+04+3.76340541E+00+1.82636932E+00+3.22499538E-02-1.22966874E-05    3
-2.55680795E-09+2.36210103E-12+2.59732915E+04+1.83256985E+01+0.00000000E+00    4
C4H71-2                 C   4H   7    0    0G   300.000  5000.000 1381.000    21
+1.07105686E+01+1.63539126E-02-5.63688038E-06+8.79591989E-10-5.12098725E-14    2
+2.21011255E+04-3.15300308E+01+1.56405993E+00+3.32162309E-02-1.59178310E-05    3
+2.92637814E-09-3.02645386E-14+2.57966120E+04+1.93052496E+01+0.00000000E+00    4
C4H71-3                 H   7C   4          G   298.150  2000.000 1000.00      1 !CWZ ADDED FROM YL CALCULATION
+4.46811308E+00+2.74302155E-02-1.21179861E-05+2.27424125E-09-1.08909321E-13    2
+1.32020300E+04+2.39088817E+00+2.79155108E-01+3.80223852E-02-1.87607474E-05    3
+5.39086588E-10+1.86579489E-12+1.43480047E+04+2.41411045E+01+0.00000000E+00    4
C4H71-3    1/13/16      C   4H   7    0    0G   300.000  5000.000 1367.000    11
+1.16977564E+01+1.53404517E-02-5.16928607E-06+7.95431212E-10-4.58914150E-14    2
+1.07395001E+04-3.82992966E+01+9.40350126E-01+3.56830321E-02-1.74384567E-05    3
+2.78964567E-09+1.78068599E-13+1.49303203E+04+2.11349333E+01+0.00000000E+00    4
C4H71-4                 H   7C   4          G   298.150  2000.000 1000.00      1 !CWZ ADDED FROM YL CALCULATION
+4.56421553E+00+2.67119686E-02-1.18632878E-05+2.28460254E-09-1.23630137E-13    2
+2.19202298E+04+4.77458878E+00+4.36415887E-01+3.87310525E-02-2.31537417E-05    3
+5.31945712E-09+2.40684882E-13+2.29703955E+04+2.58118647E+01+0.00000000E+00    4
C4H71-4                 C   4H   7    0    0G   300.000  5000.000 1389.000    21
+1.03875084E+01+1.63677264E-02-5.58416036E-06+8.65388736E-10-5.01415385E-14    2
+1.93282846E+04-2.86081068E+01+5.36903096E-01+3.66356251E-02-2.07814610E-05    3
+5.74895154E-09-6.05742821E-13+2.30645349E+04+2.53369983E+01+0.00000000E+00    4
C4H6-1                  H   6C   4          G   298.150  2000.000 1000.00      1 !CWZ ADDED FROM YL CALCULATION
+3.94365744E+00+2.61885493E-02-1.30711417E-05+3.18676492E-09-3.05127218E-13    2
+1.76368506E+04+4.59598196E+00-1.29199411E-01+4.22021279E-02-3.66747365E-05    3
+1.86446460E-08-4.10013530E-12+1.84653144E+04+2.43146241E+01+0.00000000E+00    4
SC3H5CHO                C   4H   6O   1    0G   300.000  5000.000 1396.000    21
+1.33892118E+01+1.39115420E-02-4.75820958E-06+7.38736618E-10-4.28606559E-14    2
-1.97917448E+04-4.60146004E+01+1.09372823E+00+4.43315368E-02-3.41918451E-05    3
+1.39369607E-08-2.33791460E-12-1.56745978E+04+1.94458467E+01+0.00000000E+00    4
SC3H5CO                 C   4H   5O   1    0G   300.000  5000.000 1396.000    11
+1.29925654E+01+1.22140721E-02-4.19305277E-06+6.52697685E-10-3.79407376E-14    2
-2.74782380E+03-4.51092470E+01+7.76401404E-01+4.26828436E-02-3.37881191E-05    3
+1.39128174E-08-2.33331638E-12+1.29903132E+03+1.98102013E+01+0.00000000E+00    4
AC3H5OCH2  9/ 8/14      C   4H   7O   1    0G   300.000  5000.000 1397.000    31
+1.19880368E+01+1.70263516E-02-5.78617265E-06+8.94150465E-10-5.16994613E-14    2
+3.48367473E+03-3.35860630E+01+1.20089076E+00+4.24760987E-02-2.94114641E-05    3
+1.11824860E-08-1.81309530E-12+7.26792055E+03+2.43628654E+01+0.00000000E+00    4
C4H7O2-1   9/ 8/14      C   4H   7O   1    0G   300.000  5000.000 1684.000    21
+1.12685690E+01+2.01724820E-02-7.41925667E-06+1.21275519E-09-7.30115348E-14    2
+2.13876442E+03-3.15208064E+01+5.16434924E+00+2.53427725E-02-1.39669041E-06    3
-6.00713944E-09+1.76696879E-12+5.03210693E+03+4.37441148E+00+0.00000000E+00    4
C4H7O1-4   3/30/16      C   4H   7O   1    0G   300.000  5000.000 1388.000    21
+1.33251126E+01+1.65057558E-02-5.65235890E-06+8.78319847E-10-5.09914580E-14    2
+1.91281414E+03-4.28181479E+01+2.44895430E+00+3.69423519E-02-1.77510852E-05    3
+2.64537530E-09+2.43666218E-13+6.16385921E+03+1.73174889E+01+0.00000000E+00    4
C4H7O2-1     03/16      C   4H   7O   1    0G   300.000  5000.000 1684.000    21
+1.12685690E+01+2.01724820E-02-7.41925667E-06+1.21275519E-09-7.30115348E-14    2
+2.13876442E+03-3.15208064E+01+5.16434924E+00+2.53427725E-02-1.39669041E-06    3
-6.00713944E-09+1.76696879E-12+5.03210693E+03+4.37441148E+00+0.00000000E+00    4
C4H7O2-1   9/ 8/14      C   4H   7O   1    0G   300.000  5000.000 1684.000    21
+1.12685690E+01+2.01724820E-02-7.41925667E-06+1.21275519E-09-7.30115348E-14    2
+2.13876442E+03-3.15208064E+01+5.16434924E+00+2.53427725E-02-1.39669041E-06    3
-6.00713944E-09+1.76696879E-12+5.03210693E+03+4.37441148E+00+0.00000000E+00    4
C4H7O2-1     03/16      C   4H   7O   1    0G   300.000  5000.000 1684.000    21
+1.12685690E+01+2.01724820E-02-7.41925667E-06+1.21275519E-09-7.30115348E-14    2
+2.13876442E+03-3.15208064E+01+5.16434924E+00+2.53427725E-02-1.39669041E-06    3
-6.00713944E-09+1.76696879E-12+5.03210693E+03+4.37441148E+00+0.00000000E+00    4
C4H7O2-1   9/ 8/14      C   4H   7O   1    0G   300.000  5000.000 1684.000    21
+1.12685690E+01+2.01724820E-02-7.41925667E-06+1.21275519E-09-7.30115348E-14    2
+2.13876442E+03-3.15208064E+01+5.16434924E+00+2.53427725E-02-1.39669041E-06    3
-6.00713944E-09+1.76696879E-12+5.03210693E+03+4.37441148E+00+0.00000000E+00    4
C4H7O2-1     03/16      C   4H   7O   1    0G   300.000  5000.000 1684.000    21
+1.12685690E+01+2.01724820E-02-7.41925667E-06+1.21275519E-09-7.30115348E-14    2
+2.13876442E+03-3.15208064E+01+5.16434924E+00+2.53427725E-02-1.39669041E-06    3
-6.00713944E-09+1.76696879E-12+5.03210693E+03+4.37441148E+00+0.00000000E+00    4
C4H7O2-1   9/ 8/14      C   4H   7O   1    0G   300.000  5000.000 1684.000    21
+1.12685690E+01+2.01724820E-02-7.41925667E-06+1.21275519E-09-7.30115348E-14    2
+2.13876442E+03-3.15208064E+01+5.16434924E+00+2.53427725E-02-1.39669041E-06    3
-6.00713944E-09+1.76696879E-12+5.03210693E+03+4.37441148E+00+0.00000000E+00    4
C4H7O2-1     03/16      C   4H   7O   1    0G   300.000  5000.000 1684.000    21
+1.12685690E+01+2.01724820E-02-7.41925667E-06+1.21275519E-09-7.30115348E-14    2
+2.13876442E+03-3.15208064E+01+5.16434924E+00+2.53427725E-02-1.39669041E-06    3
-6.00713944E-09+1.76696879E-12+5.03210693E+03+4.37441148E+00+0.00000000E+00    4
C4H7O2-1   9/ 8/14      C   4H   7O   1    0G   300.000  5000.000 1684.000    21
+1.12685690E+01+2.01724820E-02-7.41925667E-06+1.21275519E-09-7.30115348E-14    2
+2.13876442E+03-3.15208064E+01+5.16434924E+00+2.53427725E-02-1.39669041E-06    3
-6.00713944E-09+1.76696879E-12+5.03210693E+03+4.37441148E+00+0.00000000E+00    4
C4H7O2-1     03/16      C   4H   7O   1    0G   300.000  5000.000 1684.000    21
+1.12685690E+01+2.01724820E-02-7.41925667E-06+1.21275519E-09-7.30115348E-14    2
+2.13876442E+03-3.15208064E+01+5.16434924E+00+2.53427725E-02-1.39669041E-06    3
-6.00713944E-09+1.76696879E-12+5.03210693E+03+4.37441148E+00+0.00000000E+00    4
C4H7O2-1   9/ 8/14      C   4H   7O   1    0G   300.000  5000.000 1684.000    21
+1.12685690E+01+2.01724820E-02-7.41925667E-06+1.21275519E-09-7.30115348E-14    2
+2.13876442E+03-3.15208064E+01+5.16434924E+00+2.53427725E-02-1.39669041E-06    3
-6.00713944E-09+1.76696879E-12+5.03210693E+03+4.37441148E+00+0.00000000E+00    4
C4H7O2-1     03/16      C   4H   7O   1    0G   300.000  5000.000 1684.000    21
+1.12685690E+01+2.01724820E-02-7.41925667E-06+1.21275519E-09-7.30115348E-14    2
+2.13876442E+03-3.15208064E+01+5.16434924E+00+2.53427725E-02-1.39669041E-06    3
-6.00713944E-09+1.76696879E-12+5.03210693E+03+4.37441148E+00+0.00000000E+00    4
C4H7O2-1   9/ 8/14      C   4H   7O   1    0G   300.000  5000.000 1684.000    21
+1.12685690E+01+2.01724820E-02-7.41925667E-06+1.21275519E-09-7.30115348E-14    2
+2.13876442E+03-3.15208064E+01+5.16434924E+00+2.53427725E-02-1.39669041E-06    3
-6.00713944E-09+1.76696879E-12+5.03210693E+03+4.37441148E+00+0.00000000E+00    4
C4H7O2-1     03/16      C   4H   7O   1    0G   300.000  5000.000 1684.000    21
+1.12685690E+01+2.01724820E-02-7.41925667E-06+1.21275519E-09-7.30115348E-14    2
+2.13876442E+03-3.15208064E+01+5.16434924E+00+2.53427725E-02-1.39669041E-06    3
-6.00713944E-09+1.76696879E-12+5.03210693E+03+4.37441148E+00+0.00000000E+00    4
C4H7O2-1   9/ 8/14      C   4H   7O   1    0G   300.000  5000.000 1684.000    21
+1.12685690E+01+2.01724820E-02-7.41925667E-06+1.21275519E-09-7.30115348E-14    2
+2.13876442E+03-3.15208064E+01+5.16434924E+00+2.53427725E-02-1.39669041E-06    3
-6.00713944E-09+1.76696879E-12+5.03210693E+03+4.37441148E+00+0.00000000E+00    4
C4H7O2-1     03/16      C   4H   7O   1    0G   300.000  5000.000 1684.000    21
+1.12685690E+01+2.01724820E-02-7.41925667E-06+1.21275519E-09-7.30115348E-14    2
+2.13876442E+03-3.15208064E+01+5.16434924E+00+2.53427725E-02-1.39669041E-06    3
-6.00713944E-09+1.76696879E-12+5.03210693E+03+4.37441148E+00+0.00000000E+00    4
SC3H5OCH2-1             C   4H   7O   1    0G   300.000  5000.000 1382.000    31
+1.47022035E+01+1.55342107E-02-5.45701052E-06+8.62544885E-10-5.06734446E-14    2
+1.81294800E+03-5.05120353E+01+2.35694446E-01+4.67367652E-02-3.04880689E-05    3
+9.75216148E-09-1.23281228E-12+7.11668364E+03+2.81378517E+01+0.00000000E+00    4
C4H71-1O2  9/29/15      C   4H   7O   2    0G   300.000  5000.000 1390.000    31
+1.63738534E+01+1.62685376E-02-5.62192103E-06+8.78982520E-10-5.12510706E-14    2
-1.06318473E+03-5.69005716E+01+2.02223104E+00+4.85577506E-02-3.30293697E-05    3
+1.13406677E-08-1.57078109E-12+4.04143594E+03+2.06106646E+01+0.00000000E+00    4
C4H71-2O2  9/29/15      C   4H   7O   2    0G   300.000  5000.000 1394.000    31
+1.63565639E+01+1.61768136E-02-5.56610316E-06+8.67700997E-10-5.04886444E-14    2
-3.40245466E+03-5.75260769E+01+1.42459973E+00+5.20547601E-02-3.89440869E-05    3
+1.51726193E-08-2.42611664E-12+1.68854104E+03+2.23230947E+01+0.00000000E+00    4
C4H71-4O2  9/25/15      C   4H   7O   2    0G   300.000  5000.000 1390.000    31
+1.50240251E+01+1.72860962E-02-5.94297061E-06+9.25861430E-10-5.38461748E-14    2
+1.92460667E+02-4.85941022E+01+2.09042625E+00+4.57130080E-02-2.94815830E-05    3
+9.69604853E-09-1.30061388E-12+4.88932667E+03+2.15456077E+01+0.00000000E+00    4
C4H71-OOH4              C   4H   8O   2    0G   300.000  5000.000 1392.000    41
 1.59871304E+01 1.86028119E-02-6.40003189E-06 9.97531711E-10-5.80334203E-14    2
-1.70353450E+04-5.46227137E+01 1.31653247E+00 5.16546159E-02-3.47310922E-05    3
 1.20405755E-08-1.71650639E-12-1.17955885E+04 2.46384545E+01                   4
C4H61-3OOH4             C   4H   7O   2    0G   300.000  5000.000 1386.000    41
 1.68744844E+01 1.56488910E-02-5.46061738E-06 8.59386003E-10-5.03396686E-14    2
 7.26846315E+02-5.99891572E+01 9.87401421E-01 5.18591379E-02-3.67576063E-05    3
 1.30998708E-08-1.88471106E-12 6.32645285E+03 2.56429879E+01                   4
C4H6O1-3OOH4            C   4H   7O   3    0G   300.000  5000.000 1386.000    41
+1.95456291E+01+1.60358540E-02-5.61768950E-06+8.86341914E-10-5.20072732E-14    2
-1.12679434E+04-6.99490153E+01+3.83045773E+00+5.07388403E-02-3.42226447E-05    3
+1.13486298E-08-1.48529245E-12-5.61786232E+03+1.51509867E+01+0.00000000E+00    4
C4H6O2-1OOH4            C   4H   7O   3    0G   300.000  5000.000 1364.000    41
+2.05164800E+01+1.55727845E-02-5.54197222E-06+8.83592649E-10-5.22241946E-14    2
-9.30030707E+03-7.46630628E+01+5.38344712E+00+4.47089832E-02-2.43630482E-05    3
+5.07835349E-09-1.20805939E-13-3.40711224E+03+8.84731441E+00+0.00000000E+00    4
C4H71-3OOCH3            C   5H  10O   2    0G   300.000  5000.000 1387.000    51
+2.12299326E+01+2.07003584E-02-6.99464238E-06+1.07836941E-09-6.22999849E-14    2
-1.85005682E+04-8.53499854E+01-5.42404662E-01+7.51511469E-02-6.00684679E-05    3
+2.49701271E-08-4.22319878E-12-1.13061371E+04+3.02981962E+01+0.00000000E+00    4
C4H72-1OOCH3            C   5H  10O   2    0G   300.000  5000.000 1382.000    51
+1.92914755E+01+2.34475159E-02-8.16713690E-06+1.28338262E-09-7.50837828E-14    2
-1.72688938E+04-7.16509708E+01+2.44675386E+00+6.21430218E-02-4.39326296E-05    3
+1.72567499E-08-2.94950711E-12-1.11431755E+04+1.94028997E+01+0.00000000E+00    4
C4H8-2     8/12/15      C   4H   8    0    0G   300.000  5000.000 1383.000    21
+1.08652083E+01+1.84123129E-02-6.26886673E-06+9.70205962E-10-5.61638967E-14    2
-7.09625867E+03-3.51547481E+01+1.30795510E+00+3.53136624E-02-1.51866126E-05    3
+1.64112363E-09+3.44257620E-13-3.19767852E+03+1.81594717E+01+0.00000000E+00    4
C4H72-2                 H   7C   4          G   298.150  2000.000 1000.00      1 !CWZ ADDED 
+4.37426341E+00+2.57363050E-02-1.00546557E-05+1.27639840E-09+6.13336241E-14    2
+2.40972649E+04+4.63882080E+00+3.87261475E+00+1.94663362E-02+1.17651426E-05    3
-2.15466972E-08+7.83624839E-12+2.46114228E+04+9.12812646E+00+0.00000000E+00    4
C4H72-2    8/12/15      C   4H   7    0    0G   300.000  5000.000 1378.000    21
+1.05359634E+01+1.65535631E-02-5.71669066E-06+8.93155269E-10-5.20432637E-14    2
+2.08161211E+04-3.11046229E+01+2.46499885E+00+2.94957335E-02-1.08904521E-05    3
+9.17747264E-11+5.46417906E-13+2.42904093E+04+1.44728237E+01+0.00000000E+00    4
C4H72-2O2  9/29/15      C   4H   7O   2    0G   300.000  5000.000 1390.000    31
+1.63301022E+01+1.60698895E-02-5.50238293E-06+8.55098973E-10-4.96517196E-14    2
-4.70039715E+03-5.78736400E+01+2.49537080E+00+4.75680882E-02-3.26452548E-05    3
+1.14069694E-08-1.61494862E-12+1.76383849E+02+1.67027189E+01+0.00000000E+00    4
SC4H8OH-1               C   4H   9O   1    0G   300.000  5000.000 1405.000    41
+1.50517242E+01+1.84748629E-02-6.15327969E-06+9.38017339E-10-5.37214281E-14    2
-1.71974443E+04-5.03733848E+01+1.78282749E+00+5.18872497E-02-3.89600849E-05    3
+1.57818686E-08-2.64133852E-12-1.28305019E+04+2.00308244E+01+0.00000000E+00    4
SC4H8OH-2               C   4H   9O   1    0G   300.000  5000.000 1395.000    41
+1.45514712E+01+1.92722299E-02-6.50955109E-06+1.00200009E-09-5.77830714E-14    2
-2.09909632E+04-4.82454428E+01+1.96361387E+00+4.77673982E-02-3.11652479E-05    3
+1.07498897E-08-1.54834306E-12-1.65000330E+04+1.97286755E+01+0.00000000E+00    4
SC4H8OH-3               C   4H   9O   1    0G   300.000  5000.000 1403.000    41
+1.42453780E+01+1.89491000E-02-6.27403528E-06+9.52692609E-10-5.44157896E-14    2
-1.81803642E+04-4.56206494E+01+1.93185505E+00+4.79506224E-02-3.23719194E-05    3
+1.16232751E-08-1.72498918E-12-1.39431370E+04+2.03995003E+01+0.00000000E+00    4
SC4H8OH-1O2             C   4H   9O   3    0G   300.000  5000.000 1405.000    51
+1.88547090E+01+2.02217653E-02-6.82328766E-06+1.04961552E-09-6.05032676E-14    2
-3.65721162E+04-6.59105449E+01+1.47037864E+00+6.38295256E-02-4.92333916E-05    3
+1.99704964E-08-3.30499356E-12-3.08602292E+04+2.63462505E+01+0.00000000E+00    4
SC4H8OH-3O2             C   4H   9O   3    0G   300.000  5000.000 1417.000    51
+1.93082953E+01+1.92156764E-02-6.34250732E-06+9.60912935E-10-5.47939937E-14    2
-3.84370805E+04-6.88887622E+01+1.78918281E+00+6.62988026E-02-5.52280656E-05    3
+2.40247962E-08-4.18762027E-12-3.30428157E+04+2.28885942E+01+0.00000000E+00    4
PQC4H8OS                C   4H   9O   3    0G   300.000  5000.000 1403.000    51
+1.99993833E+01+1.96391125E-02-6.70755815E-06+1.04036085E-09-6.03187960E-14    2
-2.71257575E+04-7.31284601E+01+2.68979886E+00+6.10664073E-02-4.46910607E-05    3
+1.68939056E-08-2.59692346E-12-2.12460925E+04+1.94271757E+01+0.00000000E+00    4
PQC4H7OHS-3             C   4H   9O   3    0G   300.000  5000.000 1404.000    61
+1.89703648E+01+1.96512375E-02-6.61522830E-06+1.01590849E-09-5.84889733E-14    2
-2.92876345E+04-6.40682635E+01+3.14058820E+00+5.94343278E-02-4.55414505E-05    3
+1.85507067E-08-3.10109441E-12-2.40765022E+04+1.99412365E+01+0.00000000E+00    4
SQC4H7OHS-4             C   4H   9O   3    0G   300.000  5000.000 1414.000    61
+2.06664415E+01+1.78772156E-02-5.93193686E-06+9.02005813E-10-5.15691990E-14    2
-3.04132233E+04-7.44595459E+01+3.37952725E+00+6.50949152E-02-5.59109752E-05    3
+2.49644089E-08-4.44896795E-12-2.51501593E+04+1.58596901E+01+0.00000000E+00    4
SQC4H8OS                C   4H   9O   3    0G   300.000  5000.000 1424.000    51
+2.05363895E+01+1.85261859E-02-6.18257770E-06+9.44045247E-10-5.41390400E-14    2
-2.90453556E+04-7.66224497E+01+3.45579406E+00+6.10420456E-02-4.64106547E-05    3
+1.80687264E-08-2.81124474E-12-2.34835698E+04+1.39991890E+01+0.00000000E+00    4
NC4KET12OH              C   4H   8O   2    0G   300.000  5000.000 1384.000    41
+1.68650782E+01+1.83319076E-02-6.41389893E-06+1.01105283E-09-5.92858731E-14    2
-5.27353126E+04-5.97188408E+01+5.20269850E-01+5.40316915E-02-3.57074151E-05    3
+1.18022134E-08-1.57485744E-12-4.67781081E+04+2.89999061E+01+0.00000000E+00    4
NC4KET23OH    7/27/15   C   4H   8O   2    0G   300.000  5000.000 1386.000    41
+1.54636087E+01+1.92120108E-02-6.64681122E-06+1.03988604E-09-6.06552757E-14    2
-5.57292725E+04-5.19147488E+01+1.64761234E+00+4.74122084E-02-2.72508571E-05    3
+7.25755846E-09-6.68682869E-13-5.04946247E+04+2.37800424E+01+0.00000000E+00    4
CH3COCOHCH3             C   4H   7O   2    0G   300.000  5000.000 1395.000    41
+1.65624631E+01+1.59037217E-02-5.54554278E-06+8.72274939E-10-5.10735025E-14    2
-3.65884887E+04-6.10833920E+01-1.65607674E+00+6.08409982E-02-4.85215440E-05    3
+1.97794382E-08-3.26305133E-12-3.05158227E+04+3.58911868E+01+0.00000000E+00    4
CH3COHCO   9/24/15      C   3H   4O   2    0G   300.000  5000.000 1410.000    21
+1.50110709E+01+7.26697312E-03-2.42872486E-06+3.71246886E-10-2.13068531E-14    2
-3.87354954E+04-5.41005540E+01+8.25855205E-01+5.22217422E-02-5.66992291E-05    3
+2.94815948E-08-5.81714952E-12-3.50157127E+04+1.78488731E+01+0.00000000E+00    4
CH2COHCHO  9/24/15      C   3H   4O   2    0G   300.000  5000.000 1406.000    21
+1.40200417E+01+7.95092924E-03-2.63244516E-06+3.99896432E-10-2.28538120E-14    2
-3.76808145E+04-4.80457990E+01+5.76639663E-02+5.16589617E-02-5.49773816E-05    3
+2.83487148E-08-5.57464421E-12-3.39594513E+04+2.29757289E+01+0.00000000E+00    4
C4H71-3OH               C   4H   8O   1    0G   300.000  5000.000 1385.000    31
+1.42401634E+01+1.83038695E-02-6.37213444E-06+1.00099740E-09-5.85511411E-14    2
-2.68183960E+04-4.83949774E+01+7.16707858E-02+5.04772909E-02-3.50356983E-05    3
+1.30539199E-08-2.07783174E-12-2.16983717E+04+2.82072724E+01+0.00000000E+00    4
C4H72-2OH               C   4H   8O   1    0G   300.000  5000.000 1402.000    31
+1.49411596E+01+1.66289929E-02-5.55627511E-06+8.48898851E-10-4.86949390E-14    2
-3.12496851E+04-5.51730870E+01-1.84033728E-01+5.90104774E-02-5.22507028E-05    3
+2.44135801E-08-4.56518659E-12-2.66717960E+04+2.36075268E+01+0.00000000E+00    4
C4H63,1-3OH             C   4H   7O   1    0G   300.000  5000.000 1380.000    21
+1.33633351E+01+1.70222596E-02-5.95245190E-06+9.37896168E-10-5.49767305E-14    2
-9.90113178E+03-4.54753472E+01+5.96155469E-01+4.35893351E-02-2.65985265E-05    3
+8.14250262E-09-1.02316366E-12-5.05630797E+03+2.43923636E+01+0.00000000E+00    4
CCY(COCC)OH             C   4H   8O   2    0G   300.000  5000.000 1328.000    21
+1.03816782E+01+2.53052690E-02-1.00511826E-05+1.68204740E-09-9.58092966E-14    2
-3.94348914E+04-2.73522595E+01-6.13260697E+00+7.75376285E-02-6.73066149E-05    3
+2.82841623E-08-4.65470382E-12-3.57825027E+04+5.53089299E+01+0.00000000E+00    4
SQC4H7OHS-4O2           C   4H   9O   5    0G   300.000  5000.000 1414.000    71
+2.46607662E+01+1.92947770E-02-6.45433722E-06+9.87246207E-10-5.66889630E-14    2
-4.98467067E+04-9.10424907E+01+2.90986916E+00+7.76596028E-02-6.68513896E-05    3
+2.93627835E-08-5.12008013E-12-4.31551961E+04+2.29130715E+01+0.00000000E+00    4
C4H7O2-1,3OOH           C   4H   9O   5    0G   300.000  5000.000 1425.000    71
+2.54691227E+01+1.86441036E-02-6.23825706E-06+9.54422873E-10-5.48154425E-14    2
-4.01531561E+04-9.60389710E+01+4.88339443E+00+7.18219147E-02-5.86792171E-05    3
+2.42823866E-08-3.98538527E-12-3.36575518E+04+1.24696185E+01+0.00000000E+00    4
NC4KET13OH-2            C   4H   8O   4    0G   300.000  5000.000 1395.000    61
+2.25434165E+01+1.76377030E-02-6.14926113E-06+9.67201484E-10-5.66321794E-14    2
-6.59724022E+04-8.48522697E+01+2.13332105E+00+6.69840817E-02-5.19672275E-05    3
+2.03864253E-08-3.22074763E-12-5.90962942E+04+2.40964870E+01+0.00000000E+00    4
C4H6OHOOH1-2-3          C   4H   8O   3    0G   300.000  5000.000 1403.000    51
+2.32793098E+01+1.38280934E-02-4.61330737E-06+7.05319574E-10-4.05174739E-14    2
-4.26348237E+04-9.51979841E+01-2.88475927E+00+9.16099207E-02-9.37152074E-05    3
+4.66406895E-08-8.92736049E-12-3.52899912E+04+3.92851633E+01+0.00000000E+00    4
SC2H2OH    9/25/15      C   2H   3O   1    0G   300.000  5000.000 1410.000    11
+7.99235139E+00+5.83109353E-03-1.89242965E-06+2.83129118E-10-1.59933287E-14    2
+9.51237374E+03-1.62058375E+01+1.63791895E+00+2.64968839E-02-2.74821415E-05    3
+1.43110557E-08-2.85794966E-12+1.11467016E+04+1.58714777E+01+0.00000000E+00    4
CH2COHCO   9/25/15      C   3H   3O   2    0G   300.000  5000.000 1411.000    11
+1.31285142E+01+6.17948608E-03-1.93387986E-06+2.81892606E-10-1.56244314E-14    2
-1.93507932E+04-4.22958094E+01+1.24341370E+00+4.71484739E-02-5.44200189E-05    3
+2.95970356E-08-6.01447282E-12-1.65555219E+04+1.68301276E+01+0.00000000E+00    4
PC4H8OH-1               C   4H   9O   1    0G   300.000  5000.000 1392.000    41
+1.47813217E+01+1.89692972E-02-6.38671427E-06+9.81341181E-10-5.65332084E-14    2
-1.88487062E+04-4.98892364E+01+7.72566991E-01+5.00429367E-02-3.20163534E-05    3
+1.02913291E-08-1.30709217E-12-1.38421800E+04+2.58928300E+01+0.00000000E+00    4
PC4H8OH-2               C   4H   9O   1    0G   300.000  5000.000 1396.000    41
+1.47198620E+01+1.93691825E-02-6.59356634E-06+1.02018538E-09-5.90410746E-14    2
-1.53023402E+04-4.85296396E+01+1.89476538E+00+4.87803114E-02-3.26702980E-05    3
+1.17119949E-08-1.77100238E-12-1.07455371E+04+2.06226225E+01+0.00000000E+00    4
PC4H8OH-3               C   4H   9O   1    0G   300.000  5000.000 1398.000    41
+1.45944628E+01+1.92223378E-02-6.48868808E-06+9.98309067E-10-5.75488987E-14    2
-1.52392636E+04-4.85127747E+01+2.21685429E+00+4.71340178E-02-3.04254756E-05    3
+1.03165429E-08-1.45043599E-12-1.08208508E+04+1.83497891E+01+0.00000000E+00    4
PC4H8OH-4               C   4H   9O   1    0G   300.000  5000.000 1401.000    41
+1.41519859E+01+1.96439700E-02-6.64537615E-06+1.02402720E-09-5.91001981E-14    2
-1.56141213E+04-4.50604102E+01-6.95634735E-02+5.20263179E-02-3.44849029E-05    3
+1.17704221E-08-1.63047436E-12-1.06053581E+04+3.15909567E+01+0.00000000E+00    4
PC4H8OH-2O2             C   4H   9O   3    0G   300.000  5000.000 1407.000    51
+1.90513685E+01+2.00624257E-02-6.76970282E-06+1.04136985E-09-6.00271674E-14    2
-3.65966815E+04-6.71202048E+01+1.97780900E+00+6.25692373E-02-4.76730210E-05    3
+1.90561997E-08-3.10596799E-12-3.09625439E+04+2.35880251E+01+0.00000000E+00    4
SQC4H8OP                C   4H   9O   3    0G   300.000  5000.000 1421.000    51
+2.02482113E+01+1.90403096E-02-6.41818812E-06+9.86791658E-10-5.68666168E-14    2
-2.70686177E+04-7.43734665E+01+3.92966105E+00+5.67740736E-02-3.88077818E-05    3
+1.31554059E-08-1.72822772E-12-2.14649445E+04+1.32313419E+01+0.00000000E+00    4
SQC4H7OHP-4             C   4H   9O   3    0G   300.000  5000.000 1410.000    61
+1.99207495E+01+1.89422879E-02-6.39488327E-06+9.84231371E-10-5.67606301E-14    2
-2.89250584E+04-7.01061222E+01+1.44518283E+00+6.52944119E-02-5.10380130E-05    3
+2.05238910E-08-3.32050656E-12-2.29059890E+04+2.78546218E+01+0.00000000E+00    4
CY(CCCO)COH             C   4H   8O   2    0G   300.000  5000.000 1396.000    21
+1.34636332E+01+2.28745777E-02-9.93619553E-06+1.89605197E-09-1.26466856E-13    2
-3.96396606E+04-4.51064489E+01-6.97589766E+00+7.98392838E-02-7.11131714E-05    3
+3.16611877E-08-5.61324136E-12-3.35777839E+04+6.12093340E+01+0.00000000E+00    4
NC4KET21OH              C   4H   8O   2    0G   300.000  5000.000 1507.000    41
+1.52252911E+01+1.86615017E-02-6.30658772E-06+9.72355897E-10-5.61770184E-14    2
-5.34759661E+04-5.00397269E+01+5.46677192E+00+3.01119974E-02-2.59548850E-06    3
-7.61700554E-09+2.55573161E-12-4.89909104E+04+6.33307684E+00+0.00000000E+00    4
C2H5CHOHCO              C   4H   7O   2    0G   300.000  5000.000 1389.000    41
+1.82917246E+01+1.48007410E-02-5.24974573E-06+8.35220286E-10-4.92942253E-14    2
-3.36703722E+04-7.12363783E+01-2.44749259E+00+6.46308488E-02-5.10457937E-05    3
+1.99850773E-08-3.12214490E-12-2.66670442E+04+3.95566556E+01+0.00000000E+00    4
C2H4COCH2OH             C   4H   7O   2    0G   300.000  5000.000 1462.000    41
+1.40828195E+01+1.76833414E-02-6.09759192E-06+9.52794521E-10-5.55571628E-14    2
-3.37518398E+04-4.08944306E+01+7.98874348E+00+1.41152447E-02+1.86299924E-05    3
-1.99223089E-08+5.12983835E-12-2.98706372E+04-1.87192030E+00+0.00000000E+00    4
CH3COCHO                C   3H   4O   2    0G   300.000  5000.000 1381.000    21
+1.14371190E+01+1.06773624E-02-3.68967757E-06+5.77006752E-10-3.36532201E-14    2
-3.78079398E+04-3.25054087E+01+2.08731049E+00+3.09032484E-02-1.98794164E-05    3
+6.26174519E-09-7.69945504E-13-3.43989451E+04+1.82839639E+01+0.00000000E+00    4
C4H71-1OH               C   4H   8O   1    0G   300.000  5000.000 1402.000    31
+1.42586569E+01+1.71932504E-02-5.74956414E-06+8.79089774E-10-5.04586493E-14    2
-2.78051048E+04-4.96581579E+01-4.65981165E-01+5.56573217E-02-4.50578305E-05    3
+1.93726056E-08-3.38967639E-12-2.31007894E+04+2.79744544E+01+0.00000000E+00    4
C4H71-4OH               C   4H   8O   1    0G   300.000  5000.000 1396.000    31
+1.33437331E+01+1.82063693E-02-6.15150719E-06+9.47318576E-10-5.46543216E-14    2
-2.48479001E+04-4.27998774E+01-2.12276307E-01+4.86358034E-02-3.17241965E-05    3
+1.04986646E-08-1.39007078E-12-2.00365173E+04+3.04092052E+01+0.00000000E+00    4
C4H72-1OH               C   4H   8O   1    0G   300.000  5000.000 1367.000    31
+1.32893235E+01+1.93843938E-02-6.80733358E-06+1.07559847E-09-6.31698641E-14    2
-2.58627911E+04-4.34782359E+01+2.94637661E+00+3.45852975E-02-1.10024787E-05    3
-1.33281467E-09+9.54964043E-13-2.12241816E+04+1.55037145E+01+0.00000000E+00    4
C4H71-2OH               C   4H   8O   1    0G   300.000  5000.000 1404.000    31
+1.50658194E+01+1.65276030E-02-5.52197706E-06+8.43591643E-10-4.83870716E-14    2
-2.99737946E+04-5.53405024E+01-1.28560619E+00+6.35758020E-02-5.85328191E-05    3
+2.80452715E-08-5.32187122E-12-2.51538600E+04+2.93802791E+01+0.00000000E+00    4
C4H63,1-2OH             C   4H   7O   1    0G   300.000  5000.000 1404.000    21
+1.46899596E+01+1.48008021E-02-4.94483770E-06+7.55542892E-10-4.33461574E-14    2
-1.29448240E+04-5.45653093E+01-1.58903600E+00+6.17722944E-02-5.78263835E-05    3
+2.78090017E-08-5.26779799E-12-8.17977186E+03+2.96999338E+01+0.00000000E+00    4
C4H64,2-1OH             C   4H   7O   1    0G   300.000  5000.000 1391.000    21!CWZ UPDATES
+1.41572617E+01+1.51593460E-02-5.06194661E-06+7.74219003E-10-4.44825487E-14    2
-6.99410675E+03-4.76128315E+01-7.57727592E-01+4.98662425E-02-3.52717214E-05    3
+1.24304234E-08-1.72237947E-12-1.88378754E+03+3.24005872E+01+0.00000000E+00    4
C4H63,1-1OH             C   4H   7O   1    0G   300.000  5000.000 1401.000    21
+1.38675222E+01+1.54795810E-02-5.17720236E-06+7.91828077E-10-4.54656891E-14    2
-1.07655481E+04-4.87820652E+01-5.96640682E-01+5.31885124E-02-4.34791765E-05    3
+1.86514084E-08-3.23780972E-12-6.15543596E+03+2.74734171E+01+0.00000000E+00    4
C4H5OH-13  9/24/15      C   4H   6O   1    0G   300.000  5000.000 1405.000    21
+1.40975061E+01+1.29826578E-02-4.36356696E-06+6.69260196E-10-3.84920001E-14    2
-1.41099189E+04-4.94340793E+01-1.60022758E+00+6.12386329E-02-6.18933585E-05    3
+3.14927455E-08-6.20396658E-12-9.77435172E+03+3.08328186E+01+0.00000000E+00    4
SQC4H7OHP-4O2           C   4H   9O   5    0G   300.000  5000.000 1402.000    71
+2.35936348E+01+2.08588461E-02-7.13602285E-06+1.10820581E-09-6.43133049E-14    2
-4.78452356E+04-8.49505816E+01+2.62618431E+00+7.26812595E-02-5.64956508E-05    3
+2.25892409E-08-3.65246549E-12-4.08999596E+04+2.65615323E+01+0.00000000E+00    4
PQC4H7OHS-3O2           C   4H   9O   5    0G   300.000  5000.000 1414.000    71
+2.46607662E+01+1.92947770E-02-6.45433722E-06+9.87246207E-10-5.66889630E-14    2
-4.98467067E+04-9.10424907E+01+2.90986916E+00+7.76596028E-02-6.68513896E-05    3
+2.93627835E-08-5.12008013E-12-4.31551961E+04+2.29130715E+01+0.00000000E+00    4
NC4KET24OH-1            C   4H   8O   4    0G   300.000  5000.000 1672.000    61
+1.76639507E+01+2.38921914E-02-8.87612081E-06+1.46065294E-09-8.83476797E-14    2
-6.36561283E+04-5.60405234E+01+7.17383002E+00+3.72830917E-02-7.30000099E-06    3
-5.42423663E-09+1.94298976E-12-5.91469605E+04+3.98040888E+00+0.00000000E+00    4
NC4KET24OH-3            C   4H   8O   4    0G   300.000  5000.000 1392.000    61
+2.02237496E+01+1.94540798E-02-6.73928381E-06+1.05529414E-09-6.15931037E-14    2
-6.68651215E+04-6.99676945E+01+2.60979522E+00+6.11530456E-02-4.50409252E-05    3
+1.73313054E-08-2.75573967E-12-6.07708447E+04+2.44892030E+01+0.00000000E+00    4
C4H6OHOOH1-4-3          C   4H   8O   3    0G   300.000  5000.000 1398.000    51
+2.15163584E+01+1.55811846E-02-5.27569793E-06+8.14810620E-10-4.71424652E-14    2
-3.74825726E+04-8.24101150E+01-1.90016482E+00+7.72727339E-02-6.79667571E-05    3
+2.98158102E-08-5.16343458E-12-3.01649655E+04+4.06810164E+01+0.00000000E+00    4
C4H6OHOOH1-4-3          C   4H   8O   3    0G   300.000  5000.000 1398.000    51
+2.15163584E+01+1.55811846E-02-5.27569793E-06+8.14810620E-10-4.71424652E-14    2
-3.74825726E+04-8.24101150E+01-1.90016482E+00+7.72727339E-02-6.79667571E-05    3
+2.98158102E-08-5.16343458E-12-3.01649655E+04+4.06810164E+01+0.00000000E+00    4
C4H6OHOOH1-4-3          C   4H   8O   3    0G   300.000  5000.000 1398.000    51
+2.15163584E+01+1.55811846E-02-5.27569793E-06+8.14810620E-10-4.71424652E-14    2
-3.74825726E+04-8.24101150E+01-1.90016482E+00+7.72727339E-02-6.79667571E-05    3
+2.98158102E-08-5.16343458E-12-3.01649655E+04+4.06810164E+01+0.00000000E+00    4
C4H6OHOOH1-4-3          C   4H   8O   3    0G   300.000  5000.000 1398.000    51
+2.15163584E+01+1.55811846E-02-5.27569793E-06+8.14810620E-10-4.71424652E-14    2
-3.74825726E+04-8.24101150E+01-1.90016482E+00+7.72727339E-02-6.79667571E-05    3
+2.98158102E-08-5.16343458E-12-3.01649655E+04+4.06810164E+01+0.00000000E+00    4
C4H6OHOOH1-4-3          C   4H   8O   3    0G   300.000  5000.000 1398.000    51
+2.15163584E+01+1.55811846E-02-5.27569793E-06+8.14810620E-10-4.71424652E-14    2
-3.74825726E+04-8.24101150E+01-1.90016482E+00+7.72727339E-02-6.79667571E-05    3
+2.98158102E-08-5.16343458E-12-3.01649655E+04+4.06810164E+01+0.00000000E+00    4
C4H6OHOOH1-4-3          C   4H   8O   3    0G   300.000  5000.000 1398.000    51
+2.15163584E+01+1.55811846E-02-5.27569793E-06+8.14810620E-10-4.71424652E-14    2
-3.74825726E+04-8.24101150E+01-1.90016482E+00+7.72727339E-02-6.79667571E-05    3
+2.98158102E-08-5.16343458E-12-3.01649655E+04+4.06810164E+01+0.00000000E+00    4
C4H6OHOOH1-4-3          C   4H   8O   3    0G   300.000  5000.000 1398.000    51
+2.15163584E+01+1.55811846E-02-5.27569793E-06+8.14810620E-10-4.71424652E-14    2
-3.74825726E+04-8.24101150E+01-1.90016482E+00+7.72727339E-02-6.79667571E-05    3
+2.98158102E-08-5.16343458E-12-3.01649655E+04+4.06810164E+01+0.00000000E+00    4
C4H6OHOOH1-4-3          C   4H   8O   3    0G   300.000  5000.000 1398.000    51
+2.15163584E+01+1.55811846E-02-5.27569793E-06+8.14810620E-10-4.71424652E-14    2
-3.74825726E+04-8.24101150E+01-1.90016482E+00+7.72727339E-02-6.79667571E-05    3
+2.98158102E-08-5.16343458E-12-3.01649655E+04+4.06810164E+01+0.00000000E+00    4
C4H6OHOOH1-4-3          C   4H   8O   3    0G   300.000  5000.000 1398.000    51
+2.15163584E+01+1.55811846E-02-5.27569793E-06+8.14810620E-10-4.71424652E-14    2
-3.74825726E+04-8.24101150E+01-1.90016482E+00+7.72727339E-02-6.79667571E-05    3
+2.98158102E-08-5.16343458E-12-3.01649655E+04+4.06810164E+01+0.00000000E+00    4
C4H6OHOOH1-4-3          C   4H   8O   3    0G   300.000  5000.000 1398.000    51
+2.15163584E+01+1.55811846E-02-5.27569793E-06+8.14810620E-10-4.71424652E-14    2
-3.74825726E+04-8.24101150E+01-1.90016482E+00+7.72727339E-02-6.79667571E-05    3
+2.98158102E-08-5.16343458E-12-3.01649655E+04+4.06810164E+01+0.00000000E+00    4
C4H6OHOOH1-4-3          C   4H   8O   3    0G   300.000  5000.000 1398.000    51
+2.15163584E+01+1.55811846E-02-5.27569793E-06+8.14810620E-10-4.71424652E-14    2
-3.74825726E+04-8.24101150E+01-1.90016482E+00+7.72727339E-02-6.79667571E-05    3
+2.98158102E-08-5.16343458E-12-3.01649655E+04+4.06810164E+01+0.00000000E+00    4
C4H6OHOOH1-4-3          C   4H   8O   3    0G   300.000  5000.000 1398.000    51
+2.15163584E+01+1.55811846E-02-5.27569793E-06+8.14810620E-10-4.71424652E-14    2
-3.74825726E+04-8.24101150E+01-1.90016482E+00+7.72727339E-02-6.79667571E-05    3
+2.98158102E-08-5.16343458E-12-3.01649655E+04+4.06810164E+01+0.00000000E+00    4
C4H6OHOOH1-4-3          C   4H   8O   3    0G   300.000  5000.000 1398.000    51
+2.15163584E+01+1.55811846E-02-5.27569793E-06+8.14810620E-10-4.71424652E-14    2
-3.74825726E+04-8.24101150E+01-1.90016482E+00+7.72727339E-02-6.79667571E-05    3
+2.98158102E-08-5.16343458E-12-3.01649655E+04+4.06810164E+01+0.00000000E+00    4
C4H6OHOOH1-4-3          C   4H   8O   3    0G   300.000  5000.000 1398.000    51
+2.15163584E+01+1.55811846E-02-5.27569793E-06+8.14810620E-10-4.71424652E-14    2
-3.74825726E+04-8.24101150E+01-1.90016482E+00+7.72727339E-02-6.79667571E-05    3
+2.98158102E-08-5.16343458E-12-3.01649655E+04+4.06810164E+01+0.00000000E+00    4
C4H6OHOOH1-4-3          C   4H   8O   3    0G   300.000  5000.000 1398.000    51
+2.15163584E+01+1.55811846E-02-5.27569793E-06+8.14810620E-10-4.71424652E-14    2
-3.74825726E+04-8.24101150E+01-1.90016482E+00+7.72727339E-02-6.79667571E-05    3
+2.98158102E-08-5.16343458E-12-3.01649655E+04+4.06810164E+01+0.00000000E+00    4
C4H6OHOOH1-4-3          C   4H   8O   3    0G   300.000  5000.000 1398.000    51
+2.15163584E+01+1.55811846E-02-5.27569793E-06+8.14810620E-10-4.71424652E-14    2
-3.74825726E+04-8.24101150E+01-1.90016482E+00+7.72727339E-02-6.79667571E-05    3
+2.98158102E-08-5.16343458E-12-3.01649655E+04+4.06810164E+01+0.00000000E+00    4
C4H6OHOOH2-2-1          C   4H   8O   3    0G   300.000  5000.000 1396.000    51
+2.16656460E+01+1.59965487E-02-5.52214578E-06+8.62740322E-10-5.02768063E-14    2
-4.14875437E+04-8.39377540E+01+4.72576793E-02+7.85787048E-02-7.68006410E-05    3
+3.79206120E-08-7.33203833E-12-3.51140091E+04+2.80064858E+01+0.00000000E+00    4
C4H6OHOOH1-3-4          C   4H   8O   3    0G   300.000  5000.000 1391.000    51
+1.93445152E+01+1.82185729E-02-6.34491630E-06+9.97097673E-10-5.83420009E-14    2
-3.79952136E+04-6.88144861E+01+9.44277749E-01+6.34330602E-02-4.99455695E-05    3
+2.05720571E-08-3.48143957E-12-3.17827282E+04+2.92923796E+01+0.00000000E+00    4
HOCH2COCH2              C   3H   5O   2    0G   300.000  5000.000 1363.000    31
+1.27106963E+01+1.15513960E-02-3.95951917E-06+6.16237371E-10-3.58328248E-14    2
-2.71538154E+04-3.67129478E+01+4.98634970E+00+2.51766916E-02-1.10893306E-05    3
+1.12011467E-09+2.89491135E-13-2.40047973E+04+6.38258616E+00+0.00000000E+00    4
HOCH2CHO   9/24/15      C   2H   4O   2    0G   300.000  5000.000 1680.000    21
+7.99598542E+00+1.20664034E-02-4.43693399E-06+7.25167046E-10-4.36535460E-14    2
-4.09020567E+04-1.33754312E+01+4.35084369E+00+1.50412895E-02-5.95083030E-07    3
-3.75736217E-09+1.09353598E-12-3.91654526E+04+8.09610238E+00+0.00000000E+00    4
HOCH2CO    9/25/15      C   2H   3O   2    0G   300.000  5000.000 1487.000    21
+9.43496508E+00+7.68897340E-03-2.74959280E-06+4.39772312E-10-2.60488233E-14    2
-2.29700136E+04-2.04618579E+01+5.12916864E+00+9.07172819E-03+6.49228146E-06    3
-8.56591893E-09+2.31070825E-12-2.06151607E+04+5.73007596E+00+0.00000000E+00    4
HOCHCHO    9/25/15      C   2H   3O   2    0G   300.000  5000.000 1680.000    21
+9.99251726E+00+7.77560619E-03-2.94238616E-06+4.90136333E-10-2.98979778E-14    2
-2.20440827E+04-2.73957153E+01+5.42856274E-01+2.95295948E-02-2.08315490E-05    3
+6.72777461E-09-8.06116446E-13-1.89378452E+04+2.31681075E+01+0.00000000E+00    4
CH3COCHOH  9/25/15      C   3H   5O   2    0G   300.000  5000.000 1378.000    31
+1.23884831E+01+1.23099892E-02-4.32263800E-06+6.83043939E-10-4.01192794E-14    2
-2.97609476E+04-3.85682589E+01+2.11183979E+00+3.32521318E-02-1.96834015E-05    3
+5.40736760E-09-5.32450556E-13-2.58545486E+04+1.77643465E+01+0.00000000E+00    4
IC4H8OH-IT              C   4H   9O   1    0G   300.000  5000.000 1391.000    41
+1.29136746E+01+2.06583409E-02-6.98445966E-06+1.07562552E-09-6.20443876E-14    2
-1.81394866E+04-3.84972088E+01+3.05275715E+00+3.93926461E-02-1.90686417E-05    3
+3.86408022E-09-1.48005244E-13-1.42263749E+04+1.60840537E+01+0.00000000E+00    4
IC4H8OH-TI              C   4H   9O   1    0G   300.000  5000.000 1402.000    41
+1.46323607E+01+1.88895981E-02-6.30561450E-06+9.62474230E-10-5.51640163E-14    2
-1.87976018E+04-4.93218793E+01+2.33169342E+00+5.13017040E-02-4.02698872E-05    3
+1.75150405E-08-3.16001727E-12-1.48318978E+04+1.55368130E+01+0.00000000E+00    4
TQJC4H8OH               C   4H   9O   3    0G   300.000  5000.000 1415.000    51
+2.29681617E+01+1.65162786E-02-5.50247318E-06+8.39335285E-10-4.81030625E-14    2
-4.10051460E+04-9.34897892E+01-6.43419503E-01+8.49131517E-02-8.17210578E-05    3
+3.90979927E-08-7.27092842E-12-3.42375932E+04+2.84394025E+01+0.00000000E+00    4
TQC4H7OHI         L 2/00C   4H   9O   3    0G   300.000  5000.000 1404.000    61
+2.08281225E+01+1.81675094E-02-6.12943202E-06+9.43194119E-10-5.43937008E-14    2
-3.37386684E+04-7.74823720E+01+2.55843807E+00+6.37086077E-02-4.97169945E-05    3
+1.99225109E-08-3.21373436E-12-2.77526909E+04+1.95001368E+01+0.00000000E+00    4
IQJC4H8OH         L 2/00C   4H   9O   3    0G   300.000  5000.000 1410.000    51
+2.11752212E+01+1.75144254E-02-5.73227292E-06+8.63386596E-10-4.90282414E-14    2
-3.98881576E+04-8.19187015E+01+1.81448831E+00+7.47452750E-02-7.10895172E-05    3
+3.44973679E-08-6.54646593E-12-3.44023586E+04+1.77380434E+01+0.00000000E+00    4
TQC4H8OI                C   4H   9O   3    0G   300.000  5000.000 1411.000    51
+2.13200701E+01+1.80489663E-02-6.06124072E-06+9.29740751E-10-5.34977374E-14    2
-3.12966663E+04-8.20046659E+01+7.45747835E-02+7.46499596E-02-6.42255048E-05    3
+2.80908988E-08-4.87692045E-12-2.47182737E+04+2.94511549E+01+0.00000000E+00    4
QC4H7OHP                C   4H   9O   3    0G   300.000  5000.000 1416.000    61
+2.43481084E+01+1.50316366E-02-5.01788017E-06+7.66774357E-10-4.40093220E-14    2
-3.31922320E+04-9.68211106E+01-1.27864186E+00+8.94492926E-02-8.78565423E-05    3
+4.22110919E-08-7.83450876E-12-2.58975226E+04+3.53963909E+01+0.00000000E+00    4
IQC4H8OT                C   4H   9O   3    0G   300.000  5000.000 1405.000    51
+2.04823628E+01+1.82966721E-02-6.04413378E-06+9.16380548E-10-5.22866551E-14    2
-2.94287153E+04-7.53563247E+01+3.72211529E+00+6.42864861E-02-5.52809053E-05    3
+2.50036630E-08-4.53471908E-12-2.43110525E+04+1.21981167E+01+0.00000000E+00    4
IQC4H7OHT               C   4H   9O   3    0G   300.000  5000.000 1413.000    61
+2.19945886E+01+1.62011186E-02-5.23758492E-06+7.81898296E-10-4.41125515E-14    2
-3.07383725E+04-8.16613568E+01+3.58900054E+00+7.25591129E-02-7.14080484E-05    3
+3.55250907E-08-6.84991795E-12-2.57241250E+04+1.23766657E+01+0.00000000E+00    4
IC4H7OH                 C   4H   8O   1    0G   300.000  5000.000 1398.000    31
+1.23304221E+01+1.83885172E-02-6.06721733E-06+9.19054723E-10-5.24036171E-14    2
-2.59452023E+04-3.67418286E+01+2.04124240E+00+4.14387207E-02-2.55228632E-05    3
+8.28133017E-09-1.10654457E-12-2.22709637E+04+1.88699473E+01+0.00000000E+00    4
IC4H8OH    2/14/95 THERMC   4H   9O   1    0G   300.000  5000.000 1376.000    41
+1.25605997E+01+2.10637488E-02-7.15019648E-06+1.10439262E-09-6.38428695E-14    2
-1.86203249E+04-3.67889430E+01+3.29612707E+00+3.47649647E-02-1.02505618E-05    3
-2.04641931E-09+1.18879408E-12-1.45627247E+04+1.58606320E+01+0.00000000E+00    4
CCY(CCOC)OH       L 2/00C   4H   8O   2    0G   300.000  5000.000 1404.000    21
+1.43404718E+01+1.98311504E-02-6.60657660E-06+1.00779570E-09-5.77614335E-14    2
-4.30959414E+04-5.30535015E+01-2.84914896E+00+6.23736856E-02-4.70326536E-05    3
+1.84908286E-08-2.94976027E-12-3.74257004E+04+3.83163588E+01+0.00000000E+00    4
CCY(CCO)COH             C   4H   8O   2    0G   300.000  5000.000 1412.000    31
+1.91884885E+01+1.56255714E-02-5.22569800E-06+7.99171074E-10-4.58832445E-14    2
-4.71120302E+04-7.84579023E+01-7.10048774E+00+9.53371808E-02-9.78701612E-05    3
+4.90005646E-08-9.41685766E-12-3.98987202E+04+5.60924667E+01+0.00000000E+00    4
C2CY(COC)OH             C   4H   8O   2    0G   300.000  5000.000 1393.000    31
+1.56829970E+01+1.92910506E-02-6.63718495E-06+1.03441014E-09-6.01715267E-14    2
-4.10598236E+04-5.85686221E+01+5.92324183E-01+5.52429007E-02-4.02419018E-05    3
+1.57152217E-08-2.57388393E-12-3.58241476E+04+2.23378086E+01+0.00000000E+00    4
IC3H6OHCHO              C   4H   8O   2    0G   300.000  5000.000 1393.000    41
+1.60254376E+01+1.85402212E-02-6.36973877E-06+9.91732739E-10-5.76472640E-14    2
-5.50198923E+04-5.83074874E+01+1.84080874E+00+5.29601347E-02-3.94261774E-05    3
+1.59063430E-08-2.69565279E-12-5.01437169E+04+1.75482756E+01+0.00000000E+00    4
CH2COHCH2OOH            C   3H   6O   3    0G   300.000  5000.000 1398.000    41
+1.87971268E+01+1.12783442E-02-3.90789058E-06+6.12064651E-10-3.57305453E-14    2
-3.61154867E+04-6.94914300E+01-3.89823383E-01+7.01531131E-02-7.42036788E-05    3
+3.84181056E-08-7.63555985E-12-3.07879938E+04+2.86873505E+01+0.00000000E+00    4
TQC4H7OHIO2             C   4H   9O   5    0G   300.000  5000.000 1402.000    71
+2.82564819E+01+1.66969871E-02-5.67314614E-06+8.78350442E-10-5.09090253E-14    2
-5.66017464E+04-1.15147927E+02+3.17336206E+00+7.94005900E-02-6.51165712E-05    3
+2.62035931E-08-4.13406290E-12-4.84943162E+04+1.77867184E+01+0.00000000E+00    4
TQC4H7OHTO2             C   4H   9O   5    0G   300.000  5000.000 1402.000    71
+2.82564819E+01+1.66969871E-02-5.67314614E-06+8.78350442E-10-5.09090253E-14    2
-5.66017464E+04-1.15147927E+02+3.17336206E+00+7.94005900E-02-6.51165712E-05    3
+2.62035931E-08-4.13406290E-12-4.84943162E+04+1.77867184E+01+0.00000000E+00    4
TQC4H7OHIQ-I            C   4H   9O   5    0G   300.000  5000.000 1384.000    71
+2.88466964E+01+1.66289773E-02-5.74301906E-06+8.98791324E-10-5.24794891E-14    2
-4.69249234E+04-1.19117836E+02+6.09881562E+00+6.93745451E-02-5.12049498E-05    3
+1.81276221E-08-2.46329781E-12-3.91393707E+04+2.93862639E+00+0.00000000E+00    4
TQC4H7OHIQ-P            C   4H   9O   5    0G   300.000  5000.000 1400.000    81
+2.81439191E+01+1.63524649E-02-5.54998081E-06+8.58603978E-10-4.97359401E-14    2
-4.84502814E+04-1.11572783E+02+3.36947511E+00+7.96855226E-02-6.74365765E-05    3
+2.82233283E-08-4.65270820E-12-4.05567534E+04+1.92726029E+01+0.00000000E+00    4
IQC4H7OHTO2             C   4H   9O   5    0G   300.000  5000.000 1389.000    71
+2.41720261E+01+2.09397176E-02-7.29061406E-06+1.14554056E-09-6.70217517E-14    2
-5.04772118E+04-8.95996685E+01+3.83287364E+00+6.90926177E-02-5.15031144E-05    3
+1.99235553E-08-3.17456897E-12-4.34442789E+04+1.94648622E+01+0.00000000E+00    4
IQC4H8OTQ-I             C   4H   9O   5    0G   300.000  5000.000 1386.000    71
+2.53249383E+01+2.00634820E-02-7.01249558E-06+1.10475030E-09-6.47561724E-14    2
-4.09610593E+04-9.73592779E+01+5.90219800E+00+6.26952142E-02-4.17351838E-05    3
+1.35422162E-08-1.71169663E-12-3.39620020E+04+7.89290087E+00+0.00000000E+00    4
IQC4H7OHTQ-P            C   4H   9O   5    0G   300.000  5000.000 1391.000    81
+2.45769593E+01+2.01889393E-02-7.03584537E-06+1.10623327E-09-6.47523225E-14    2
-4.25783112E+04-9.05052742E+01+3.45242802E+00+7.14541224E-02-5.54616790E-05    3
+2.22754676E-08-3.66067450E-12-3.54133076E+04+2.23024492E+01+0.00000000E+00    4
CH2CQCOHQ  7/ 1/14      C   3H   6O   5    0G   300.000  5000.000 1418.000    61
+3.86574091E+01+4.83815026E-04-2.10413843E-07+3.81490832E-11-2.46187754E-15    2
-6.56392184E+04-1.61083579E+02-1.61171759E+01+1.78866440E-01-2.16751308E-04    3
+1.15450289E-07-2.27163078E-11-5.21165145E+04+1.14441286E+02+0.00000000E+00    4
IC3H5COHQ               C   4H   8O   3    0G   300.000  5000.000 1504.000    51
+2.07387831E+01+1.58360934E-02-5.27614462E-06+8.05932218E-10-4.62682425E-14    2
-4.41821241E+04-7.94239893E+01+2.64360992E+00+5.72485066E-02-3.95907807E-05    3
+1.27775635E-08-1.47241476E-12-3.80099993E+04+1.77322273E+01+0.00000000E+00    4
IC3H5Q                  C   3H   6O   2    0G   300.000  5000.000 1397.000    31
+1.43424294E+01+1.28053632E-02-4.40584813E-06+6.86848148E-10-3.99675209E-14    2
-1.65261025E+04-4.89934539E+01+1.32903007E+00+4.49170722E-02-3.51235127E-05    3
+1.41982181E-08-2.33335008E-12-1.21898396E+04+2.02696565E+01+0.00000000E+00    4
COHQCYC(COC)            C   4H   8O   4    0G   300.000  5000.000 1319.000    51
+2.44599226E+01+1.64187782E-02-5.74024372E-06+9.05710407E-10-5.31829152E-14    2
-6.01811228E+04-1.02049722E+02+2.40687943E+00+5.95180442E-02-3.16913659E-05    3
+4.23694824E-09+8.42033474E-13-5.19694864E+04+1.88941416E+01+0.00000000E+00    4
QCYC(CCOC)OH            C   4H   8O   4    0G   300.000  5000.000 1411.000    41
+2.20860197E+01+1.83743733E-02-6.29478769E-06+9.78787994E-10-5.68621317E-14    2
-5.89652037E+04-8.64964494E+01-2.09099972E+00+8.02656739E-02-6.69756245E-05    3
+2.79282034E-08-4.60981823E-12-5.12529252E+04+4.11897260E+01+0.00000000E+00    4
HOCOCQ(CH3)2            C   4H   8O   4    0G   300.000  5000.000 1380.000    61
+2.28935401E+01+1.78627606E-02-6.34627520E-06+1.01068546E-09-5.96885712E-14    2
-8.05400680E+04-9.08953779E+01+1.56326363E+00+6.77165643E-02-5.14600149E-05    3
+1.99184629E-08-3.16007445E-12-7.30943302E+04+2.37255421E+01+0.00000000E+00    4
CHOC(CH3)OHCH2Q         C   4H   8O   4    0G   300.000  5000.000 1383.000    61
+2.24480753E+01+1.78753902E-02-6.26904597E-06+9.90084046E-10-5.81417382E-14    2
-6.55093075E+04-8.56747327E+01+2.40933530E+00+6.13326038E-02-4.03874986E-05    3
+1.22738404E-08-1.32997480E-12-5.83049516E+04+2.29870742E+01+0.00000000E+00    4
CO(CH2OOH)2             C   3H   6O   5    0G   300.000  5000.000 1393.000    61
+2.43376341E+01+1.14074110E-02-4.08931881E-06+6.55183244E-10-3.88570518E-14    2
-5.16862647E+04-9.01518175E+01-2.47626577E+00+8.93736793E-02-9.25891121E-05    3
+4.63168490E-08-8.93300309E-12-4.38924057E+04+4.84479477E+01+0.00000000E+00    4
C4H6                    H   6C   4          G   298.150  2000.000 1000.00      1 !CWZ ADDED FROM YL CALCULATION
+6.48731037E+00+2.20209540E-02-9.83379092E-06+1.91675967E-09-1.06427710E-13    2
+1.01596660E+04-1.06711837E+01-3.37272121E+00+5.76700106E-02-5.76207712E-05    3
+2.99836767E-08-6.17538953E-12+1.23212258E+04+3.78455365E+01+0.00000000E+00    4
C4H5-I                  H  5 C  4 O  0      G     298.0    3000.0    1000.0    1
 5.25595308E+00 2.19965949E-02-1.09137173E-05 2.63404317E-09-2.50557472E-13    2
 3.57055213E+04-1.56386290E+00-4.20623364E-01 4.38861302E-02-4.32708486E-05    3
 2.43849315E-08-5.85727339E-12 3.69066616E+04 2.60889512E+01                   4
C4H5-N                  H  5 C  4 O  0      G     298.0    3000.0    1000.0    1
 7.29521441E+00 1.91513156E-02-9.57154022E-06 2.33661465E-09-2.25148097E-13    2
 4.01314083E+04-1.35255263E+01-3.18360247E+00 5.81813715E-02-6.38641527E-05    3
 3.57450182E-08-7.89217819E-12 4.23740398E+04 3.77564497E+01                   4
C3H3CH2OOH   12/16      C   4H   6O   2    0G   300.000  5000.000 1384.000    31
 1.76337943E+01 1.27580284E-02-4.44136954E-06 6.98375539E-10-4.08987084E-14    2
 4.20746041E+03-6.27097953E+01 1.64825356E+00 5.28806082E-02-4.39833841E-05    3
 1.88140805E-08-3.26453253E-12 9.50410156E+03 2.21988630E+01                   4
C3H3CH2O  10/12/16      C   4H   5O   1    0G   300.000  5000.000 1676.000    11
 1.14427994E+01 1.50893347E-02-5.59321856E-06 9.19032913E-10-5.55290838E-14    2
 2.35239513E+04-3.19110047E+01 5.53696698E+00 2.18274562E-02-3.15173599E-06    3
-3.93256542E-09 1.28730350E-12 2.61457576E+04 2.17741565E+00                   4
C3H3CHO   10/12/16      C   4H   4O   1    0G   300.000  5000.000 1395.000    11
 1.27526772E+01 1.00631883E-02-3.49308972E-06 5.47746784E-10-3.20020827E-14    2
 1.41528612E+03-4.14481197E+01 1.14170208E+00 4.05129134E-02-3.49445730E-05    3
 1.55825190E-08-2.79824627E-12 5.13366022E+03 1.97621650E+01                   4
CYHEXDN13  8/31/16      C   6H   8    0    0G   300.000  5000.000 1392.000    01
 1.50997866E+01 2.12080269E-02-7.33544206E-06 1.14760359E-09-6.69433814E-14    2
 4.44900608E+03-6.16788333E+01-4.82039387E+00 6.70223856E-02-4.73487895E-05    3
 1.69645503E-08-2.45944445E-12 1.14209741E+04 4.55310016E+01                   4
CYHEXDN14  8/31/16      C   6H   8    0    0G   300.000  5000.000 1385.000    01
 1.57263000E+01 2.09982638E-02-7.33474543E-06 1.15498418E-09-6.76769598E-14    2
 4.37984609E+03-6.64317549E+01-3.02043825E+00 6.10388887E-02-3.86837660E-05    3
 1.17505763E-08-1.35178604E-12 1.12646687E+04 3.55809099E+01                   4
C6H8       8/31/16      C   6H   8    0    0G   300.000  5000.000 1397.000    21
 1.69511085E+01 1.86092892E-02-6.39483993E-06 9.95781471E-10-5.78882385E-14    2
 1.19358759E+04-6.63328076E+01-2.80216545E+00 7.45728595E-02-6.92665672E-05    3
 3.34618343E-08-6.42278211E-12 1.79188255E+04 3.64469277E+01                   4
CYHEXEN-4J 8/31/16      C   6H   9    0    0G   300.000  5000.000 1388.000    01
 1.45726981E+01 2.41687737E-02-8.34933859E-06 1.30512039E-09-7.60857953E-14    2
 1.40406544E+04-5.59995158E+01-3.84381292E+00 5.99346158E-02-3.11377445E-05    3
 5.82015177E-09 8.64222393E-14 2.11060274E+04 4.53885355E+01                   4
CYPENTN-4MJ             C   6H   9    0    0G10.000    3000.000  433.34        1 !W.GREEN'S
-2.41048175E+00 6.21591818E-02-3.89684972E-05 1.17648713E-08-1.36838719E-12    2 !W.GREEN'S
 2.57204512E+04 3.77632099E+01 3.94469866E+00 3.44171538E-03 1.64472094E-04    3 !W.GREEN'S
-3.01509598E-07 1.79533574E-10 2.51701784E+04 1.24235238E+01                   4 !W.GREEN'S
CYPENTN-4M4J            C   6H   9    0    0G10.000    3000.000  528.91        1 !W.GREEN'S
-3.37191907E+00 6.18953322E-02-3.77368199E-05 1.10138910E-08-1.23709218E-12    2 !W.GREEN'S
 2.17495406E+04 4.18567684E+01 4.00036055E+00-6.25727801E-04 1.58764283E-04    3 !W.GREEN'S
-2.60854825E-07 1.38700145E-10 2.10643320E+04 1.18801829E+01                   4 !W.GREEN'S
CYPENTN-4M3J            C   6H   9    0    0G10.000    3000.000  451.07        1 !W.GREEN'S
-3.01888829E+00 6.53666245E-02-4.25401593E-05 1.32583714E-08-1.58143371E-12    2 !W.GREEN'S
 1.74262118E+04 3.99119184E+01 3.94632666E+00 3.28517048E-03 1.64955619E-04    3 !W.GREEN'S
-2.94963183E-07 1.70105404E-10 1.68010595E+04 1.18895739E+01                   4 !W.GREEN'S
CYPENTN-4MTHNE          C   6H   8    0    0G10.000    3000.000  592.29        1 !W.GREEN'S
-2.10239098E+00 5.81365770E-02-3.60082225E-05 1.06656333E-08-1.21248223E-12    2 !W.GREEN'S
 1.53559396E+04 3.49539705E+01 4.03826412E+00-4.04316353E-03 1.73911296E-04    3 !W.GREEN'S
-2.84646912E-07 1.48353104E-10 1.49917771E+04 1.16115412E+01                   4 !W.GREEN'S
C4H5-2            H6W/94C   4H   5    0    0G   300.000  5000.000 1385.000    11
+1.03230828E+01+1.17625574E-02-4.00004665E-06+6.18727929E-10-3.58083530E-14    2
+3.25861413E+04-2.88794317E+01+2.31011292E+00+2.83747046E-02-1.63836755E-05    3
+4.46251967E-09-4.30510879E-13+3.55842945E+04+1.49105965E+01+0.00000000E+00    4
C4H4              H6W/94C   4H   4    0    0G   300.000  3000.00  1000.00      1
+6.65070920E+00+1.61294340E-02-7.19388750E-06+1.49817870E-09-1.18641100E-13    2
+3.11959920E+04-9.79521180E+00-1.91524790E+00+5.27508780E-02-7.16559440E-05    3
+5.50724230E-08-1.72862280E-11+3.29785040E+04+3.14199830E+01+0.00000000E+00    4
C4H3-I            AB1/93C   4H   3    0    0G   300.000  3000.00  1000.00      1
+9.09781650E+00+9.22071190E-03-3.38784410E-06+4.91604980E-10-1.45297800E-14    2
+5.66005740E+04-1.98025970E+01+2.08304120E+00+4.08342740E-02-6.21596850E-05    3
+5.16793580E-08-1.70291840E-11+5.80051290E+04+1.36174620E+01+0.00000000E+00    4
C4H3-N            H6W/94C   4H   3    0    0G   300.000  3000.00  1000.00      1
+5.43282790E+00+1.68609810E-02-9.43131090E-06+2.57038950E-09-2.74563090E-13    2
+6.16006800E+04-1.56739810E+00-3.16841130E-01+4.69121000E-02-6.80938100E-05    3
+5.31799210E-08-1.65230050E-11+6.24761990E+04+2.46225590E+01+0.00000000E+00    4
C4H2              D11/99C   4H   2    0    0G   300.000  3000.000 1000.        1
+9.15763280E+00+5.54305180E-03-1.35916040E-06+1.87800750E-11+2.31895360E-14    2
+5.25880390E+04-2.37114600E+01+1.05439780E+00+4.16269600E-02-6.58717840E-05    3
+5.32570750E-08-1.66831620E-11+5.41852110E+04+1.48665910E+01+0.00000000E+00    4
CHCC(CH2)CHCH2  16      C   6H   6    0    0G   300.000  5000.000 1386.000    21
+1.50259784E+01+1.56363629E-02-5.48046599E-06+8.64876878E-10-5.07521932E-14    2
+3.26003690E+04-5.46018534E+01-9.74937292E-02+5.25465475E-02-4.13131445E-05    3
+1.72824473E-08-3.00750335E-12+3.77892668E+04+2.62208973E+01+0.00000000E+00    4
CH2CHCHCHCCH 03/16      C   6H   6    0    0G   300.000  5000.000 1394.000    21
+1.71155812E+01+1.35873582E-02-4.71347534E-06+7.38927269E-10-4.31678854E-14    2
+3.34001333E+04-6.63949871E+01-1.63758241E+00+6.58049292E-02-6.19478129E-05    3
+2.95388753E-08-5.56039075E-12+3.91068149E+04+3.13986448E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1385.000    11
+1.39299886E+01+1.13228814E-02-3.87393567E-06+6.02378620E-10-3.50120301E-14    2
-2.39589898E+03-4.79026849E+01+4.51553480E-01+4.37530418E-02-3.37273602E-05    3
+1.31111496E-08-2.04732021E-12+2.14943141E+03+2.40835867E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1385.000    11
+1.39299886E+01+1.13228814E-02-3.87393567E-06+6.02378620E-10-3.50120301E-14    2
-2.39589898E+03-4.79026849E+01+4.51553480E-01+4.37530418E-02-3.37273602E-05    3
+1.31111496E-08-2.04732021E-12+2.14943141E+03+2.40835867E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1385.000    11
+1.39299886E+01+1.13228814E-02-3.87393567E-06+6.02378620E-10-3.50120301E-14    2
-2.39589898E+03-4.79026849E+01+4.51553480E-01+4.37530418E-02-3.37273602E-05    3
+1.31111496E-08-2.04732021E-12+2.14943141E+03+2.40835867E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1385.000    11
+1.39299886E+01+1.13228814E-02-3.87393567E-06+6.02378620E-10-3.50120301E-14    2
-2.39589898E+03-4.79026849E+01+4.51553480E-01+4.37530418E-02-3.37273602E-05    3
+1.31111496E-08-2.04732021E-12+2.14943141E+03+2.40835867E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1385.000    11
+1.39299886E+01+1.13228814E-02-3.87393567E-06+6.02378620E-10-3.50120301E-14    2
-2.39589898E+03-4.79026849E+01+4.51553480E-01+4.37530418E-02-3.37273602E-05    3
+1.31111496E-08-2.04732021E-12+2.14943141E+03+2.40835867E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1385.000    11
+1.39299886E+01+1.13228814E-02-3.87393567E-06+6.02378620E-10-3.50120301E-14    2
-2.39589898E+03-4.79026849E+01+4.51553480E-01+4.37530418E-02-3.37273602E-05    3
+1.31111496E-08-2.04732021E-12+2.14943141E+03+2.40835867E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1385.000    11
+1.39299886E+01+1.13228814E-02-3.87393567E-06+6.02378620E-10-3.50120301E-14    2
-2.39589898E+03-4.79026849E+01+4.51553480E-01+4.37530418E-02-3.37273602E-05    3
+1.31111496E-08-2.04732021E-12+2.14943141E+03+2.40835867E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1385.000    11
+1.39299886E+01+1.13228814E-02-3.87393567E-06+6.02378620E-10-3.50120301E-14    2
-2.39589898E+03-4.79026849E+01+4.51553480E-01+4.37530418E-02-3.37273602E-05    3
+1.31111496E-08-2.04732021E-12+2.14943141E+03+2.40835867E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1385.000    11
+1.39299886E+01+1.13228814E-02-3.87393567E-06+6.02378620E-10-3.50120301E-14    2
-2.39589898E+03-4.79026849E+01+4.51553480E-01+4.37530418E-02-3.37273602E-05    3
+1.31111496E-08-2.04732021E-12+2.14943141E+03+2.40835867E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1385.000    11
+1.39299886E+01+1.13228814E-02-3.87393567E-06+6.02378620E-10-3.50120301E-14    2
-2.39589898E+03-4.79026849E+01+4.51553480E-01+4.37530418E-02-3.37273602E-05    3
+1.31111496E-08-2.04732021E-12+2.14943141E+03+2.40835867E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1385.000    11
+1.39299886E+01+1.13228814E-02-3.87393567E-06+6.02378620E-10-3.50120301E-14    2
-2.39589898E+03-4.79026849E+01+4.51553480E-01+4.37530418E-02-3.37273602E-05    3
+1.31111496E-08-2.04732021E-12+2.14943141E+03+2.40835867E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1385.000    11
+1.39299886E+01+1.13228814E-02-3.87393567E-06+6.02378620E-10-3.50120301E-14    2
-2.39589898E+03-4.79026849E+01+4.51553480E-01+4.37530418E-02-3.37273602E-05    3
+1.31111496E-08-2.04732021E-12+2.14943141E+03+2.40835867E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1385.000    11
+1.39299886E+01+1.13228814E-02-3.87393567E-06+6.02378620E-10-3.50120301E-14    2
-2.39589898E+03-4.79026849E+01+4.51553480E-01+4.37530418E-02-3.37273602E-05    3
+1.31111496E-08-2.04732021E-12+2.14943141E+03+2.40835867E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1385.000    11
+1.39299886E+01+1.13228814E-02-3.87393567E-06+6.02378620E-10-3.50120301E-14    2
-2.39589898E+03-4.79026849E+01+4.51553480E-01+4.37530418E-02-3.37273602E-05    3
+1.31111496E-08-2.04732021E-12+2.14943141E+03+2.40835867E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1385.000    11
+1.39299886E+01+1.13228814E-02-3.87393567E-06+6.02378620E-10-3.50120301E-14    2
-2.39589898E+03-4.79026849E+01+4.51553480E-01+4.37530418E-02-3.37273602E-05    3
+1.31111496E-08-2.04732021E-12+2.14943141E+03+2.40835867E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1385.000    11
+1.39299886E+01+1.13228814E-02-3.87393567E-06+6.02378620E-10-3.50120301E-14    2
-2.39589898E+03-4.79026849E+01+4.51553480E-01+4.37530418E-02-3.37273602E-05    3
+1.31111496E-08-2.04732021E-12+2.14943141E+03+2.40835867E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1385.000    11
+1.39299886E+01+1.13228814E-02-3.87393567E-06+6.02378620E-10-3.50120301E-14    2
-2.39589898E+03-4.79026849E+01+4.51553480E-01+4.37530418E-02-3.37273602E-05    3
+1.31111496E-08-2.04732021E-12+2.14943141E+03+2.40835867E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1385.000    11
+1.39299886E+01+1.13228814E-02-3.87393567E-06+6.02378620E-10-3.50120301E-14    2
-2.39589898E+03-4.79026849E+01+4.51553480E-01+4.37530418E-02-3.37273602E-05    3
+1.31111496E-08-2.04732021E-12+2.14943141E+03+2.40835867E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1385.000    11
+1.39299886E+01+1.13228814E-02-3.87393567E-06+6.02378620E-10-3.50120301E-14    2
-2.39589898E+03-4.79026849E+01+4.51553480E-01+4.37530418E-02-3.37273602E-05    3
+1.31111496E-08-2.04732021E-12+2.14943141E+03+2.40835867E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1385.000    11
+1.39299886E+01+1.13228814E-02-3.87393567E-06+6.02378620E-10-3.50120301E-14    2
-2.39589898E+03-4.79026849E+01+4.51553480E-01+4.37530418E-02-3.37273602E-05    3
+1.31111496E-08-2.04732021E-12+2.14943141E+03+2.40835867E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1385.000    11
+1.39299886E+01+1.13228814E-02-3.87393567E-06+6.02378620E-10-3.50120301E-14    2
-2.39589898E+03-4.79026849E+01+4.51553480E-01+4.37530418E-02-3.37273602E-05    3
+1.31111496E-08-2.04732021E-12+2.14943141E+03+2.40835867E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1385.000    11
+1.39299886E+01+1.13228814E-02-3.87393567E-06+6.02378620E-10-3.50120301E-14    2
-2.39589898E+03-4.79026849E+01+4.51553480E-01+4.37530418E-02-3.37273602E-05    3
+1.31111496E-08-2.04732021E-12+2.14943141E+03+2.40835867E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1385.000    11
+1.39299886E+01+1.13228814E-02-3.87393567E-06+6.02378620E-10-3.50120301E-14    2
-2.39589898E+03-4.79026849E+01+4.51553480E-01+4.37530418E-02-3.37273602E-05    3
+1.31111496E-08-2.04732021E-12+2.14943141E+03+2.40835867E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1385.000    11
+1.39299886E+01+1.13228814E-02-3.87393567E-06+6.02378620E-10-3.50120301E-14    2
-2.39589898E+03-4.79026849E+01+4.51553480E-01+4.37530418E-02-3.37273602E-05    3
+1.31111496E-08-2.04732021E-12+2.14943141E+03+2.40835867E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1385.000    11
+1.39299886E+01+1.13228814E-02-3.87393567E-06+6.02378620E-10-3.50120301E-14    2
-2.39589898E+03-4.79026849E+01+4.51553480E-01+4.37530418E-02-3.37273602E-05    3
+1.31111496E-08-2.04732021E-12+2.14943141E+03+2.40835867E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1385.000    11
+1.39299886E+01+1.13228814E-02-3.87393567E-06+6.02378620E-10-3.50120301E-14    2
-2.39589898E+03-4.79026849E+01+4.51553480E-01+4.37530418E-02-3.37273602E-05    3
+1.31111496E-08-2.04732021E-12+2.14943141E+03+2.40835867E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1400.000    11
+1.32551859E+01+1.19066619E-02-4.06547591E-06+6.30312610E-10-3.65301442E-14    2
+4.28822305E+03-4.47690775E+01-4.93209912E-01+5.26550104E-02-5.15159642E-05    3
+2.57409661E-08-5.03442115E-12+8.26367547E+03+2.61133171E+01+0.00000000E+00    4
CH2CHCHCHO              C   4H   5O   1    0G   300.000  5000.000 1385.000    11
+1.39299886E+01+1.13228814E-02-3.87393567E-06+6.02378620E-10-3.50120301E-14    2
-2.39589898E+03-4.79026849E+01+4.51553480E-01+4.37530418E-02-3.37273602E-05    3
+1.31111496E-08-2.04732021E-12+2.14943141E+03+2.40835867E+01+0.00000000E+00    4
NC4H5O2                 C   4H   5O   2    0G   300.000  5000.000 1396.000    21
+1.64522106E+01+1.16956821E-02-4.08000295E-06+6.41912007E-10-3.75906771E-14    2
+1.25380689E+04-5.87190920E+01+6.12413489E-01+5.52512502E-02-5.12447815E-05    3
+2.41307414E-08-4.50077091E-12+1.74115237E+04+2.40736828E+01+0.00000000E+00    4
C2H3CHOHCH2             C   4H   7O   1    0G   300.000  5000.000 1382.000    31
+1.44787895E+01+1.56397705E-02-5.47239981E-06+8.62563884E-10-5.05719495E-14    2
-1.47613624E+03-4.69553537E+01+2.30466478E+00+4.41216304E-02-3.23935804E-05    3
+1.31499701E-08-2.29928167E-12+2.89743860E+03+1.86657957E+01+0.00000000E+00    4
C2H3CHOHCH2OO           C   4H   7O   3    0G   300.000  5000.000 1389.000    41
+1.83530129E+01+1.69514703E-02-5.91054392E-06+9.29544125E-10-5.44175546E-14    2
-2.07620807E+04-6.33248942E+01+1.85132718E+00+5.68751205E-02-4.37973133E-05    3
+1.77010151E-08-2.95624741E-12-1.51170708E+04+2.48996326E+01+0.00000000E+00    4
C4H6OH1-4OOH 10/16      C   4H   8O   3    0G   300.000  5000.000 1391.000    51
 1.93445152E+01 1.82185729E-02-6.34491630E-06 9.97097673E-10-5.83420009E-14    2
-3.79952136E+04-6.88144861E+01 9.44277749E-01 6.34330602E-02-4.99455695E-05    3
 2.05720571E-08-3.48143957E-12-3.17827282E+04 2.92923796E+01                   4
C4H5OH1-4OOH 10/16      C   4H   7O   3    0G   300.000  5000.000 1388.000    51
 1.91838037E+01 1.59285036E-02-5.58251870E-06 8.81016733E-10-5.17029398E-14    2
-1.00934916E+04-6.62734801E+01 2.30965628E+00 5.66530089E-02-4.39894466E-05    3
 1.77261106E-08-2.93544265E-12-4.32625775E+03 2.39530949E+01                   4
C4H6OH1-2,4OOH 10/16    C   4H   8O   5    0G   300.000  5000.000 1394.000    71
 2.57425089E+01 1.72396246E-02-6.05608891E-06 9.57322306E-10-5.62477620E-14    2
-5.28215509E+04-9.80930757E+01 1.50567086E+00 8.08823060E-02-7.14931886E-05    3
 3.19609885E-08-5.69861501E-12-4.51133784E+04 2.95736160E+01                   4
C4H5OH1-4OOH-2OO        C   4H   7O   5    0G   300.000  5000.000 1393.000    61
 2.47662773E+01 1.59483622E-02-5.61098009E-06 8.87848597E-10-5.22018160E-14    2
-3.55928552E+04-9.19981196E+01 2.31183130E+00 7.47918419E-02-6.60490378E-05    3
 2.95219734E-08-5.26743325E-12-2.84330075E+04 2.63334617E+01                   4
C4H5OH1-2,4OOH 10/16    C   4H   7O   5    0G   300.000  5000.000 1389.000    71
 2.37938036E+01 1.63846860E-02-5.76911110E-06 9.13313993E-10-5.37158479E-14    2
-2.98477456E+04-8.42153079E+01 3.64255921E+00 6.68210812E-02-5.52639509E-05    3
 2.34596615E-08-4.03883583E-12-2.31592732E+04 2.28638284E+01                   4
C4H5OJ1-2,4OOH 10/16    C   4H   7O   5    0G   300.000  5000.000 1392.000    61
 2.59610037E+01 1.50317787E-02-5.31796267E-06 8.44637677E-10-4.97916701E-14    2
-2.60964572E+04-9.93170329E+01 4.33801022E+00 6.85025374E-02-5.62798005E-05    3
 2.30600805E-08-3.77375439E-12-1.89425384E+04 1.56651703E+01                   4
C3H3OHCHO1-2OOH         C   4H   6O   4    0G   300.000  5000.000 1671.000    51
 2.01194396E+01 1.68368880E-02-6.36172689E-06 1.05867042E-09-6.45335884E-14    2
-4.78792303E+04-7.27686560E+01 1.79127621E+00 5.72787740E-02-3.75143238E-05    3
 1.08389158E-08-1.07752428E-12-4.16873725E+04 2.59257566E+01                   4
C3H4CH2OH-3O            C   4H   7O   2    0G   300.000  5000.000 1384.000    31
+1.67237902E+01+1.62893097E-02-5.69978133E-06+8.98524197E-10-5.26886310E-14    2
-1.90975797E+04-5.73256364E+01+2.45139062E+00+4.76173501E-02-3.17417435E-05    3
+1.07287265E-08-1.48712660E-12-1.38958927E+04+2.01150648E+01+0.00000000E+00    4
C2H3CHOHCH2OOH          C   4H   8O   3    0G   300.000  5000.000 1391.000    51
 1.93445152E+01 1.82185729E-02-6.34491630E-06 9.97097673E-10-5.83420009E-14    2
-3.79952136E+04-6.88144861E+01 9.44277749E-01 6.34330602E-02-4.99455695E-05    3
 2.05720571E-08-3.48143957E-12-3.17827282E+04 2.92923796E+01                   4
C4H51,3OH2  ENOL  T12/15C  4.H  6.O  1.   0.G   200.000  6000.000 1000.        1
 1.17568770E+01 1.62957646E-02-5.86745770E-06 9.47794368E-10-5.68012244E-14    2
-1.33808588E+04-3.61322949E+01 5.32202847E-01 3.47944440E-02 9.07363332E-06    3
-4.26890292E-08 2.13649260E-11-9.76102764E+03 2.46259582E+01-8.04995700E+03    4
C2H3CHOHCHO   9/16      C   4H   6O   2    0G   300.000  5000.000 1519.000    31
 1.62609725E+01 1.46912093E-02-5.27966798E-06 8.47240068E-10-5.03008110E-14    2
-3.45597776E+04-5.86214663E+01 1.98300140E+00 3.57502763E-02-8.68562950E-06    3
-5.68946121E-09 2.40246806E-12-2.84547220E+04 2.22890748E+01                   4
C3H3OH    11/ 9/16      C   3H   4O   1    0G   300.000  5000.000 1409.000    11
 1.07170529E+01 8.56985387E-03-2.82907434E-06 4.28605740E-10-2.44382142E-14    2
-1.98468165E+03-3.12883184E+01 6.64863235E-01 3.90790884E-02-3.85723070E-05    3
 1.92354298E-08-3.72429095E-12 8.00157434E+02 2.01988440E+01                   4
CDY(COCC)OH   9/16      C   4H   6O   2    0G   300.000  5000.000 1404.000    11
 1.59912606E+01 1.48926281E-02-5.14765273E-06 8.05057203E-10-4.69530524E-14    2
-2.64939381E+04-5.94930361E+01-4.28737799E+00 6.85313676E-02-6.01513042E-05    3
 2.65620353E-08-4.65128316E-12-2.01441601E+04 4.70823318E+01                   4
C3H2OHCH2Q    9/16      C   4H   6O   3    0G   300.000  5000.000 1386.000    41
 1.81132272E+01 1.45656351E-02-5.07825128E-06 7.98650178E-10-4.67560629E-14    2
-1.76332305E+04-6.30842082E+01 4.69903114E+00 4.54113058E-02-3.24594006E-05    3
 1.20345879E-08-1.84997432E-12-1.28888049E+04 9.19557638E+00                   4
C2H3CHOHCH2OH 9/16      C   4H   8O   2    0G   300.000  5000.000 1392.000    41
 1.63773228E+01 1.84895764E-02-6.40907987E-06 1.00394106E-09-5.86083740E-14    2
-4.57454068E+04-5.53052098E+01-2.78850131E-01 5.91275862E-02-4.54587885E-05    3
 1.85462925E-08-3.13811396E-12-4.00697341E+04 3.36435671E+01                   4
C2H3CHOHCH2O  9/16      C   4H   7O   2    0G   300.000  5000.000 1384.000    31
 1.67237902E+01 1.62893097E-02-5.69978133E-06 8.98524197E-10-5.26886310E-14    2
-1.90975797E+04-5.73256364E+01 2.45139062E+00 4.76173501E-02-3.17417435E-05    3
 1.07287265E-08-1.48712660E-12-1.38958927E+04 2.01150648E+01                   4
C2H3COCH2Q    7/16      C   4H   6O   3    0G   300.000  5000.000 1390.000    41
 2.03130199E+01 1.30620215E-02-4.64429563E-06 7.40055113E-10-4.37242482E-14    2
-3.20078211E+04-7.53059526E+01-1.68971987E+00 7.27107744E-02-6.82564997E-05    3
 3.19924185E-08-5.91996843E-12-2.51697616E+04 3.99766836E+01                   4
C3H4OCH2OH              C   4H   7O   2    0G   300.000  5000.000 1678.000    31
+1.35768442E+01+1.93824171E-02-6.93534320E-06+1.11509393E-09-6.64283563E-14    2
-2.37032565E+04-4.05883301E+01+3.68556748E+00+3.71954683E-02-1.57927917E-05    3
+1.29414603E-09+4.50053262E-13-1.99630755E+04+1.41318611E+01+0.00000000E+00    4
C2H3OCHCH2OH            C   4H   7O   2    0G   300.000  5000.000 1406.000    41
+1.61335254E+01+1.57030233E-02-5.34935592E-06+8.28273404E-10-4.79651847E-14    2
-1.69967975E+04-5.26511117E+01-2.35771595E+00+6.64956454E-02-5.97594106E-05    3
+2.74521100E-08-5.00266740E-12-1.13587733E+04+4.39223977E+01+0.00000000E+00    4
CH2CH2COCH2OH           C   4H   7O   2    0G   300.000  5000.000 1498.000    41
+1.45572634E+01+1.67757761E-02-5.67488345E-06+8.75536866E-10-5.06066052E-14    2
-2.83118087E+04-4.36209150E+01+5.86369173E+00+2.65549901E-02-1.46596470E-06    3
-7.41455041E-09+2.42515138E-12-2.42760164E+04+6.74620320E+00+0.00000000E+00    4
C2H3COCH2OH             C   4H   6O   2    0G   300.000  5000.000 1374.000    31
+1.45010066E+01+1.57293771E-02-5.52878496E-06+8.74135857E-10-5.13615582E-14    2
-3.95492218E+04-4.65251707E+01+3.52503727E+00+3.70498105E-02-2.04866837E-05    3
+5.38095100E-09-5.47927324E-13-3.51894190E+04+1.41521904E+01+0.00000000E+00    4
C3H4CH2OH-1OOH          C   4H   8O   3    0G   300.000  5000.000 1373.000    51
+2.05562405E+01+1.73434658E-02-6.08615888E-06+9.61896332E-10-5.65238760E-14    2
-3.61100647E+04-7.48563094E+01+2.62447134E+00+5.66513196E-02-3.85852510E-05    3
+1.31139830E-08-1.80853978E-12-2.95875423E+04+2.24313053E+01+0.00000000E+00    4
C3H4CH2OH-1O            C   4H   7O   2    0G   300.000  5000.000 1502.000    31
+1.71974002E+01+1.64461405E-02-5.88477087E-06+9.41603116E-10-5.57896598E-14    2
-1.83089012E+04-6.07872595E+01+6.65239296E+00+2.39519793E-02+8.12599943E-06    3
-1.51386006E-08+4.29644312E-12-1.29560218E+04+1.89176185E+00+0.00000000E+00    4
CH2OC3H4OH              C   4H   7O   2    0G   300.000  5000.000 1380.000    31
+1.55246652E+01+1.72695515E-02-6.02881277E-06+9.48883834E-10-5.55788127E-14    2
-1.61651202E+04-4.92916169E+01+2.88677533E+00+4.28670375E-02-2.48859484E-05    3
+6.91428514E-09-7.31772975E-13-1.13113370E+04+2.00967837E+01+0.00000000E+00    4
CHOC3H4OH               C   4H   6O   2    0G   300.000  5000.000 1380.000    31
+1.56483679E+01+1.46897907E-02-5.15632446E-06+8.14600326E-10-4.78399746E-14    2
-3.88944658E+04-5.34469355E+01+2.11996229E+00+4.43238416E-02-2.97127304E-05    3
+1.00484103E-08-1.39027193E-12-3.39592163E+04+1.99769992E+01+0.00000000E+00    4
C4H71-OO3               C   4H   7O   2    0G   300.000  5000.000 1391.000    31
+1.82801163E+01+1.42612723E-02-4.85633823E-06+7.52827804E-10-4.36658356E-14    2
-1.26079889E+03-6.93661163E+01-6.97499481E-01+6.24502522E-02-5.21064763E-05    3
+2.19339967E-08-3.68635153E-12+4.87666022E+03+3.10773529E+01+0.00000000E+00    4
C4H61-OOH34     16      C   4H   8O   4    0G   300.000  5000.000 1394.000    61
 2.43681963E+01 1.56262504E-02-5.36622026E-06 8.36672539E-10-4.87261234E-14    2
-2.97395130E+04-9.53858126E+01-5.50389828E-01 8.08980233E-02-7.14917402E-05    3
 3.14214570E-08-5.45705442E-12-2.18931780E+04 3.57719063E+01                   4
C4H61-OOH3-OO4  16      C   4H   7O   4    0G   300.000  5000.000 1393.000    51
 2.33277335E+01 1.44238222E-02-4.95806165E-06 7.73525973E-10-4.50682556E-14    2
-1.24821576E+04-8.89214747E+01 2.83626299E-01 7.47135230E-02-6.59702203E-05    3
 2.89687939E-08-5.02779526E-12-5.21758836E+03 3.23977640E+01                   4
C4H61-2OOH34    16      C   4H   7O   4    0G   300.000  5000.000 1392.000    61
 2.40461895E+01 1.35992427E-02-4.71882979E-06 7.40795046E-10-4.33461797E-14    2
-1.77729681E+03-9.19448524E+01 8.07371622E-01 7.42390637E-02-6.59005046E-05    3
 2.89287584E-08-5.01113774E-12 5.56275422E+03 3.04532122E+01                   4
C4H6-OOH234     16      C   4H   8O   6    0G   300.000  5000.000 1398.000    81
 3.06605815E+01 1.48149843E-02-5.14984670E-06 8.09528022E-10-4.74147104E-14    2
-4.45213885E+04-1.24066059E+02-9.72395895E-02 9.89577364E-02-9.41326054E-05    3
 4.35896844E-08-7.86256542E-12-3.52104814E+04 3.65299347E+01                   4
C4H61-OOH34-OO2 16      C   4H   7O   6    0G   300.000  5000.000 1397.000    71
 2.96189216E+01 1.36224652E-02-4.74693365E-06 7.47380161E-10-4.38219621E-14    2
-2.72652141E+04-1.17599351E+02 7.32401155E-01 9.27972124E-02-8.86481619E-05    3
 4.11651984E-08-7.44082707E-12-1.85343774E+04 3.31749869E+01                   4
C4H412-OOH34    16      C   4H   6O   4    0G   300.000  5000.000 1390.000    51
 2.37714316E+01 1.22691980E-02-4.37585634E-06 6.98707223E-10-4.13399756E-14    2
-1.05419085E+04-9.05795816E+01 2.25296705E+00 7.03405671E-02-6.59546939E-05    3
 3.07772261E-08-5.66772762E-12-3.83724444E+03 2.22442095E+01                   4
C3H3CHO-OOH23   16      C   4H   6O   5    0G   300.000  5000.000 1387.000    61
 2.70408781E+01 1.19361788E-02-4.33840618E-06 7.01448748E-10-4.18636928E-14    2
-4.19006207E+04-1.07701779E+02 1.21286535E+00 7.32715332E-02-5.85847446E-05    3
 2.18420551E-08-3.09398790E-12-3.32531372E+04 3.02888053E+01                   4
C4H4O-OOH24     16      C   4H   6O   5    0G   300.000  5000.000 1388.000    61
 2.52105579E+01 1.33311572E-02-4.78042241E-06 7.66051638E-10-4.54376448E-14    2
-3.85672545E+04-9.41153859E+01 9.59575596E-01 7.65313711E-02-6.90784876E-05    3
 3.08837168E-08-5.46998241E-12-3.08308409E+04 3.37582000E+01                   4
C4H61-4OOH3             C   4H   7O   2    0G   300.000  5000.000 1393.000    41
+1.88083591E+01+1.34574643E-02-4.59376133E-06+7.13321256E-10-4.14238605E-14    2
+6.59898017E+03-7.01085955E+01-5.85215644E-01+6.35552472E-02-5.46196793E-05    3
+2.35377539E-08-4.02918330E-12+1.27800498E+04+3.22244808E+01+0.00000000E+00    4
C4H512-OO4   03/16 THERMC   4H   5O   2    0G   300.000  5000.000 1400.000    21
+1.42836297E+01+1.30646729E-02-4.44620310E-06+6.87917196E-10-3.98144345E-14    2
+2.10779108E+04-4.44989804E+01+1.52191421E+00+4.71698948E-02-4.03200254E-05    3
+1.80912888E-08-3.27484097E-12+2.50993362E+04+2.25474610E+01+0.00000000E+00    4
CH2CCO                  H   2C   3O   1     G   298.150  2000.000 1000.00      1
 4.40003435E+00 1.25785246E-02-5.91887918E-06 1.27758857E-09-9.45874595E-14    2
 1.33314103E+04 4.29517065E+00 3.60551892E+00 1.45152309E-02-6.96190546E-06    3
 7.31583992E-10 3.52252542E-13 1.35523812E+04 8.43858717E+00                   4
C4H62-OOH14     16      C   4H   8O   4    0G   300.000  5000.000 1383.000    61
 2.40027956E+01 1.69211626E-02-6.02147599E-06 9.59977296E-10-5.67352934E-14    2
-2.74866767E+04-9.09248026E+01 5.33887384E-01 7.75331204E-02-6.82132680E-05    3
 3.07798871E-08-5.60160434E-12-1.98197385E+04 3.32306388E+01                   4
C4H513-OO2   03/16 THERMC   4H   5O   2    0G   300.000  5000.000 1405.000    21
+1.56904837E+01+1.19260796E-02-4.06874172E-06+6.30816230E-10-3.65702642E-14    2
+1.32535118E+04-5.61395385E+01-7.53229326E-01+5.71867156E-02-5.24258034E-05    3
+2.41573152E-08-4.38383698E-12+1.82311643E+04+2.96637047E+01+0.00000000E+00    4
CYCCCOO-3J   03/16 THERMC   4H   5O   2    0G   300.000  5000.000 1403.000    01
+1.47511170E+01+1.36105988E-02-4.65772901E-06+7.23551244E-10-4.20014564E-14    2
+9.03032818E+03-5.37988385E+01-2.47556740E+00+6.02141116E-02-5.37658895E-05    3
+2.43859766E-08-4.38845640E-12+1.43437053E+04+3.64073667E+01+0.00000000E+00    4
CH2CYCOO-CH2 03/16 THERMC   4H   5O   2    0G   300.000  5000.000 1398.000    21
+1.58989765E+01+1.20316212E-02-4.16546349E-06+6.52021319E-10-3.80466500E-14    2
+1.80307061E+04-5.73648764E+01+2.58755552E-01+5.57836767E-02-5.23131171E-05    3
+2.49455274E-08-4.69840113E-12+2.27704741E+04+2.41236108E+01+0.00000000E+00    4
C2H3COOCH2   03/16 THERMC   4H   5O   2    0G   300.000  5000.000 1378.000    31
+1.65803208E+01+1.15439736E-02-4.11631882E-06+6.57144442E-10-3.88749935E-14    2
-2.11309534E+04-6.07009305E+01+2.00791111E+00+4.51755954E-02-3.38733412E-05    3
+1.27342296E-08-1.94378047E-12-1.60205295E+04+1.77255740E+01+0.00000000E+00    4
CYCOOC-CH2   03/16 THERMC   4H   5O   2    0G   300.000  5000.000 1403.000    11
+1.49632112E+01+1.28724587E-02-4.37191522E-06+6.75553099E-10-3.90654123E-14    2
+2.28933543E+04-5.25926129E+01-2.66210588E-01+5.57788088E-02-5.16416215E-05    3
+2.44394027E-08-4.56852993E-12+2.74516568E+04+2.66023034E+01+0.00000000E+00    4
C4H6O25           T 3/97C   4H   6O   1    0G   200.000  5000.000  1000.0      1
+8.60658242E+00+2.08310051E-02-8.42229481E-06+1.56717640E-09-1.09391202E-13    2
-1.76177415E+04-2.32464750E+01+2.67053463E+00+4.92586420E-03+8.86967406E-05    3
-1.26219194E-07+5.23991321E-11-1.46572472E+04+1.45722395E+01-1.30831522E+04    4
C2H3CHOCH2              C   4H   6O   1    0G   300.000  5000.000 1431.000    11
+1.26762790E+01+1.40819509E-02-4.63473868E-06+7.01090838E-10-3.99438277E-14    2
-4.08065264E+03-4.22515995E+01-3.59388437E+00+5.79063450E-02-4.97163294E-05    3
+2.15818682E-08-3.69199072E-12+8.58852628E+02+4.28475443E+01+0.00000000E+00    4
C4H4O             T03/97C   4H   4O   1    0G   200.000  6000.0    1000.0      1
+9.38935003E+00+1.40291241E-02-5.07755110E-06+8.24137332E-10-4.95319963E-14    2
-8.68241814E+03-2.79162920E+01+8.47469463E-01+1.31773796E-02+5.99735901E-05    3
-9.71562904E-08+4.22733796E-11-5.36785445E+03+2.14945172E+01-4.17166616E+03    4
C4H6O23           T 3/97C   4H   6O   1    0G   200.000  5000.000  1000.0      1
+8.60658242E+00+2.08310051E-02-8.42229481E-06+1.56717640E-09-1.09391202E-13    2
-1.32392815E+04-2.32464750E+01+2.67053463E+00+4.92586420E-03+8.86967406E-05    3
-1.26219194E-07+5.23991321E-11-1.02787872E+04+1.45722395E+01-1.30831522E+04    4
C4H612                  H   6C   4          G   298.150  2000.000 1000.00      1 !CWZ ADDED FROM YL CALCULATION
+4.03554835E+00+2.50965369E-02-1.14318520E-05+2.30461618E-09-1.42764873E-13    2
+1.69864966E+04+4.60107412E+00+1.26299208E+00+3.21839229E-02-1.60586721E-05    3
+1.38632371E-09+1.08751804E-12+1.77411498E+04+1.89777653E+01+0.00000000E+00    4
C4H612            A 8/83C   4H   6    0    0G   300.000  5000.000 1374.000    11
+1.14059885E+01+1.31489843E-02-4.43542071E-06+6.83028825E-10-3.94289265E-14    2
+1.42427294E+04-3.69674067E+01+9.45515689E-01+3.46162239E-02-1.98590697E-05    3
+5.02139421E-09-3.67977164E-13+1.81439079E+04+2.02191143E+01+0.00000000E+00    4
C4H6-2                  H   6C   4          G   298.150  2000.000 1000.00      1 !CWZ ADDED FROM YL CALCULATION
+3.28493310E+00+2.56208578E-02-1.13437876E-05+2.13794807E-09-1.05016221E-13    2
+1.53435097E+04+7.73047992E+00+2.65653419E+00+2.30439838E-02+1.57227991E-07    3
-1.06198653E-08+4.35705454E-12+1.57237129E+04+1.20347588E+01+0.00000000E+00    4
C4H6-2            A 8/83C   4H   6    0    0G   300.000  5000.000 1377.000    21
+9.60305554E+00+1.48972169E-02-5.16751230E-06+8.09757170E-10-4.72817668E-14    2
+1.24831314E+04-2.87129792E+01+1.97152408E+00+2.76790997E-02-1.13396645E-05    3
+1.02970745E-09+2.75290944E-13+1.57283766E+04+1.42147356E+01+0.00000000E+00    4
H2C4O             120189H   2C   4O   1     G  0300.00   4000.00  1000.00      1
+1.02688800E+01+4.89616400E-03-4.88508100E-07-2.70856600E-10+5.10701300E-14    2
+2.34690300E+04-2.81598500E+01+4.81097100E+00+1.31399900E-02+9.86507300E-07    3
-6.12072000E-09+1.64000300E-12+2.54580300E+04+2.11342400E+00+0.00000000E+00    4
NC3H7CHO   8/12/15      C   4H   8O   1    0G   300.000  5000.000 1679.000    31
+1.19789345E+01+2.04894148E-02-7.24831619E-06+1.15561709E-09-6.84119824E-14    2
-3.09272130E+04-3.63929716E+01+1.24208539E+00+4.21277518E-02-2.13832135E-05    3
+4.22614614E-09-1.03710908E-13-2.71049353E+04+2.21567167E+01+0.00000000E+00    4
NC3H7CO                 C   4H   7O   1    0G   300.000  5000.000 1496.000    31
+1.34870098E+01+1.58626861E-02-5.41698905E-06+8.40508889E-10-4.87570090E-14    2
-1.30725285E+04-4.38634081E+01+2.63537828E+00+3.40368642E-02-1.24118988E-05    3
-1.17886666E-09+1.16488136E-12-8.65919992E+03+1.68407569E+01+0.00000000E+00    4
C3H6CHO-1               C   4H   7O   1    0G   300.000  5000.000 1538.000    31
+1.33449137E+01+1.59347421E-02-5.43143577E-06+8.41706117E-10-4.87847084E-14    2
-6.91281947E+03-4.19662475E+01+2.21483383E+00+3.54113290E-02-1.44082892E-05    3
+5.27605922E-11+8.95003230E-13-2.46482792E+03+2.00076022E+01+0.00000000E+00    4
C3H6CHO-2               C   4H   7O   1    0G   300.000  5000.000 1439.000    31
+1.27128605E+01+1.68632757E-02-5.83779932E-06+9.14059755E-10-5.33575736E-14    2
-8.50165835E+03-3.84620358E+01+4.01372834E+00+2.33173718E-02+5.72463585E-06    3
-1.27182841E-08+3.69912722E-12-4.16766399E+03+1.30545921E+01+0.00000000E+00    4
C3H6CHO-3               C   4H   7O   1    0G   300.000  5000.000 1678.000    31
+1.21729663E+01+1.80056550E-02-6.43783092E-06+1.03362049E-09-6.14850407E-14    2
-1.08642352E+04-3.80322250E+01+5.29001237E-01+4.30707499E-02-2.49474118E-05    3
+6.40934608E-09-5.27769846E-13-6.87667117E+03+2.48856420E+01+0.00000000E+00    4
C2H5COCH3  8/12/15      C   4H   8O   1    0G   300.000  5000.000 1454.000    31
+1.28183044E+01+1.79874386E-02-5.94194784E-06+9.01636365E-10-5.14993729E-14    2
-3.51711964E+04-4.11609193E+01+2.57048052E+00+3.51446793E-02-1.23849584E-05    3
-1.21280927E-09+1.16163555E-12-3.10194049E+04+1.61395232E+01+0.00000000E+00    4
C2H5COCH2               C   4H   7O   1    0G   300.000  5000.000 1396.000    31
+1.35979480E+01+1.57187785E-02-5.35200820E-06+8.28428039E-10-4.79645862E-14    2
-1.30111973E+04-4.46215708E+01+1.96643032E+00+4.10271409E-02-2.56193885E-05    3
+7.86244495E-09-9.26825962E-13-8.80149212E+03+1.84803948E+01+0.00000000E+00    4
CH2CH2COCH3             C   4H   7O   1    0G   300.000  5000.000 1392.000    31
+1.17915603E+01+1.70296457E-02-5.75444256E-06+8.86035114E-10-5.11070778E-14    2
-9.70683178E+03-3.25532787E+01+2.36191763E+00+3.50400641E-02-1.70487065E-05    3
+3.09070210E-09+2.80364847E-14-6.02754073E+03+1.95184512E+01+0.00000000E+00    4
CH3CHCOCH3              C   4H   7O   1    0G   300.000  5000.000 1438.000    31
+1.19651378E+01+1.63142163E-02-5.39879520E-06+8.20454677E-10-4.69197541E-14    2
-1.51990676E+04-3.30142593E+01+3.31082456E+00+2.83712402E-02-5.64603859E-06    3
-4.62626296E-09+1.82954207E-12-1.14602301E+04+1.62217415E+01+0.00000000E+00    4
C2H3COCH3               C   4H   6O   1    0G   300.000  5000.000 1390.000    21
+1.19989844E+01+1.52616304E-02-5.26018882E-06+8.20774274E-10-4.77834528E-14    2
-2.12170620E+04-3.71383523E+01+6.55910700E-01+4.19405303E-02-3.00269693E-05    3
+1.16578089E-08-1.92100897E-12-1.72216627E+04+2.38412293E+01+0.00000000E+00    4
CH3CHOOCOCH3            C   4H   7O   3    0G   300.000  5000.000 1411.000    41
+1.68056216E+01+1.70791389E-02-5.69439450E-06+8.68878944E-10-4.98008338E-14    2
-3.06718613E+04-5.51178960E+01+4.30171569E+00+4.62273591E-02-3.12564494E-05    3
+1.08627824E-08-1.51478379E-12-2.63732146E+04+1.19724375E+01+0.00000000E+00    4
CH2CHOOHCOCH3           C   4H   7O   3    0G   300.000  5000.000 1413.000    51
+1.78031394E+01+1.60286227E-02-5.38152372E-06+8.25242310E-10-4.74718968E-14    2
-2.30767899E+04-5.87370258E+01+4.45962223E+00+4.67200276E-02-3.15878907E-05    3
+1.06245787E-08-1.38857032E-12-1.84720686E+04+1.29655977E+01+0.00000000E+00    4
C2H5CHCO                C   4H   6O   1    0G   300.000  5000.000 1550.000    21
-2.04040652E+02+2.93466880E-01-1.15884523E-04+1.95253673E-08-1.19030791E-12    2
+8.27380036E+04+1.21233386E+03-2.28307043E+01+1.70978191E-01-3.53394379E-04    3
+2.78221616E-07-6.77325074E-11-1.04125457E+04+1.31232921E+02+0.00000000E+00    4
NC5H12     9/ 8/14      C   5H  12    0    0G   300.000  5000.000 1393.000    41
+1.58289132E+01+2.59344752E-02-8.83016276E-06+1.36654986E-09-7.91029283E-14    2
-2.59397429E+04-6.05558457E+01-2.99551806E-01+5.94963054E-02-3.41764359E-05    3
+9.47896058E-09-9.73675086E-13-1.98959978E+04+2.75742132E+01+0.00000000E+00    4
C5H11-1    9/ 8/14      C   5H  11    0    0G   300.000  5000.000 1394.000    41
+1.51918481E+01+2.40339049E-02-8.19717624E-06+1.27002751E-09-7.35727956E-14    2
-8.02148517E+02-5.36479311E+01+9.83190194E-02+5.58653605E-02-3.28855625E-05    3
+9.58366873E-09-1.08641370E-12+4.82065818E+03+2.86921367E+01+0.00000000E+00    4
C5H11-2    9/ 8/14      C   5H  11    0    0G   300.000  5000.000 1395.000    41
+1.47177050E+01+2.41667557E-02-8.18647646E-06+1.26271867E-09-7.29267957E-14    2
-2.26027771E+03-5.06071115E+01+8.17689455E-01+4.92653514E-02-2.13785619E-05    3
+1.85532454E-09+7.06259101E-13+3.26221492E+03+2.65876082E+01+0.00000000E+00    4
C5H11-3    9/ 8/14      C   5H  11    0    0G   300.000  5000.000 1395.000    41
+1.47177050E+01+2.41667557E-02-8.18647646E-06+1.26271867E-09-7.29267957E-14    2
-2.26027771E+03-5.12965931E+01+8.17689455E-01+4.92653514E-02-2.13785619E-05    3
+1.85532454E-09+7.06259101E-13+3.26221492E+03+2.58981266E+01+0.00000000E+00    4
C5H11O2H-1 9/ 8/14      C   5H  12O   2    0G   300.000  5000.000 1393.000    61
+2.08826791E+01+2.61587380E-02-8.96860003E-06+1.39463023E-09-8.10033260E-14    2
-3.71864314E+04-8.01917306E+01+7.56966700E-01+7.13994143E-02-4.75006334E-05    3
+1.62337006E-08-2.26834390E-12-3.00009521E+04+2.85558826E+01+0.00000000E+00    4
C5H11O2H-2 9/ 8/14      C   5H  12O   2    0G   300.000  5000.000 1400.000    61
+2.11347974E+01+2.56494323E-02-8.72650240E-06+1.34983451E-09-7.81086942E-14    2
-3.90416300E+04-8.21964012E+01+1.06841342E+00+7.36472213E-02-5.31234084E-05    3
+2.02380955E-08-3.18671855E-12-3.21746715E+04+2.51901593E+01+0.00000000E+00    4
C5H11O2H-3 9/ 8/14      C   5H  12O   2    0G   300.000  5000.000 1400.000    61
+2.11347974E+01+2.56494323E-02-8.72650240E-06+1.34983451E-09-7.81086942E-14    2
-3.90416300E+04-8.35753644E+01+1.06841342E+00+7.36472213E-02-5.31234084E-05    3
+2.02380955E-08-3.18671855E-12-3.21746715E+04+2.38111961E+01+0.00000000E+00    4
C5H11O2-1  9/ 8/14      C   5H  11O   2    0G   300.000  5000.000 1392.000    51
+1.99508904E+01+2.48182054E-02-8.50415197E-06+1.32191009E-09-7.67596518E-14    2
-1.99782879E+04-7.43587406E+01+1.47849612E+00+6.56222617E-02-4.24002295E-05    3
+1.39455731E-08-1.86035665E-12-1.33065245E+04+2.57184992E+01+0.00000000E+00    4
C5H11O2-2  9/ 8/14      C   5H  11O   2    0G   300.000  5000.000 1401.000    51
+2.01379084E+01+2.43048677E-02-8.24744582E-06+1.27344965E-09-7.35953601E-14    2
-2.17777897E+04-7.59194124E+01+1.95945265E+00+6.73012650E-02-4.74261817E-05    3
+1.76453313E-08-2.71599328E-12-1.55102022E+04+2.15326067E+01+0.00000000E+00    4
C5H11O2-3  9/ 8/14      C   5H  11O   2    0G   300.000  5000.000 1401.000    51
+2.01379084E+01+2.43048677E-02-8.24744582E-06+1.27344965E-09-7.35953601E-14    2
-2.17777897E+04-7.72983757E+01+1.95945265E+00+6.73012650E-02-4.74261817E-05    3
+1.76453313E-08-2.71599328E-12-1.55102022E+04+2.01536434E+01+0.00000000E+00    4
C5H11O-1   9/ 8/14      C   5H  11O   1    0G   300.000  5000.000 1396.000    41
+1.87118024E+01+2.36054696E-02-8.05610528E-06+1.24900841E-09-7.23989034E-14    2
-1.84133036E+04-7.11769229E+01+1.61443159E+00+5.84449099E-02-3.26027513E-05    3
+7.76525028E-09-4.48739932E-13-1.20210227E+04+2.23620687E+01+0.00000000E+00    4
C5H11O-2   9/ 8/14      C   5H  11O   1    0G   300.000  5000.000 1407.000    41
+1.85178187E+01+2.33560329E-02-7.87896503E-06+1.21190761E-09-6.98572825E-14    2
-2.01488741E+04-7.05224357E+01+1.80797841E+00+5.95687062E-02-3.62936785E-05    3
+1.05785660E-08-1.11086649E-12-1.41294991E+04+2.01085450E+01+0.00000000E+00    4
C5H11O-3   9/ 8/14      C   5H  11O   1    0G   300.000  5000.000 1407.000    41
+1.85178187E+01+2.33560329E-02-7.87896503E-06+1.21190761E-09-6.98572825E-14    2
-2.01488741E+04-7.19013990E+01+1.80797841E+00+5.95687062E-02-3.62936785E-05    3
+1.05785660E-08-1.11086649E-12-1.41294991E+04+1.87295817E+01+0.00000000E+00    4
C5H10OOH1-2 9/8/14      C   5H  11O   2    0G   300.000  5000.000 1396.000    61
+2.00795991E+01+2.43589475E-02-8.36202795E-06+1.30140406E-09-7.56329790E-14    2
-1.33166011E+04-7.30604965E+01+2.65531081E+00+6.13777489E-02-3.72526890E-05    3
+1.10683497E-08-1.26575773E-12-6.87569412E+03+2.18610512E+01+0.00000000E+00    4
C5H10OOH1-3 9/8/14      C   5H  11O   2    0G   300.000  5000.000 1396.000    61
+1.94584083E+01+2.46031733E-02-8.38534822E-06+1.29883762E-09-7.52367289E-14    2
-1.33548974E+04-6.90616123E+01+2.21641946E+00+5.96426514E-02-3.30151174E-05    3
+7.82801873E-09-4.53626906E-13-6.89038067E+03+2.53165655E+01+0.00000000E+00    4
C5H10OOH1-4 9/8/14      C   5H  11O   2    0G   300.000  5000.000 1396.000    61
+1.94584083E+01+2.46031733E-02-8.38534822E-06+1.29883762E-09-7.52367289E-14    2
-1.33548974E+04-6.90616123E+01+2.21641946E+00+5.96426514E-02-3.30151174E-05    3
+7.82801873E-09-4.53626906E-13-6.89038067E+03+2.53165655E+01+0.00000000E+00    4
C5H10OOH1-5 9/8/14      C   5H  11O   2    0G   300.000  5000.000 1393.000    61
+2.02627427E+01+2.43041392E-02-8.36491479E-06+1.30408546E-09-7.58781596E-14    2
-1.20792388E+04-7.41332935E+01+9.60306204E-01+6.85338215E-02-4.72580697E-05    3
+1.69913164E-08-2.53055987E-12-5.25227210E+03+2.99005842E+01+0.00000000E+00    4
C5H10OOH2-1 9/8/14      C   5H  11O   2    0G   300.000  5000.000 1401.000    61
+2.11683533E+01+2.30995637E-02-7.85421525E-06+1.21454488E-09-7.02697376E-14    2
-1.41652579E+04-7.96524097E+01+1.97482622E+00+6.85026751E-02-4.88793184E-05    3
+1.80505063E-08-2.71515676E-12-7.58936343E+03+2.31709703E+01+0.00000000E+00    4
C5H10OOH2-3 9/8/14      C   5H  11O   2    0G   300.000  5000.000 1410.000    61
+2.03599510E+01+2.36444020E-02-8.00996599E-06+1.23543694E-09-7.13457143E-14    2
-1.51264004E+04-7.50912668E+01+3.03844851E+00+6.35523371E-02-4.29455468E-05    3
+1.50665567E-08-2.16139351E-12-9.06691319E+03+1.81118164E+01+0.00000000E+00    4
C5H10OOH2-4 9/8/14      C   5H  11O   2    0G   300.000  5000.000 1410.000    61
+1.98843630E+01+2.37470675E-02-7.98273943E-06+1.22497373E-09-7.04946509E-14    2
-1.52413050E+04-7.19593692E+01+2.69411113E+00+6.13272504E-02-3.77802938E-05    3
+1.11809673E-08-1.20043769E-12-9.09500363E+03+2.11388648E+01+0.00000000E+00    4
C5H10OOH2-5 9/8/14      C   5H  11O   2    0G   300.000  5000.000 1401.000    61
+2.05595155E+01+2.35923560E-02-8.01736916E-06+1.23918525E-09-7.16674070E-14    2
-1.39059417E+04-7.62751847E+01+1.46239008E+00+7.00773603E-02-5.18935110E-05    3
+2.03023923E-08-3.27212476E-12-7.45896384E+03+2.56255897E+01+0.00000000E+00    4
C5H10OOH3-1 9/8/14      C   5H  11O   2    0G   300.000  5000.000 1401.000    61
+2.05595155E+01+2.35923560E-02-8.01736916E-06+1.23918525E-09-7.16674070E-14    2
-1.39059417E+04-7.69646663E+01+1.46239008E+00+7.00773603E-02-5.18935110E-05    3
+2.03023923E-08-3.27212476E-12-7.45896384E+03+2.49361080E+01+0.00000000E+00    4
C5H10OOH3-2 9/8/14      C   5H  11O   2    0G   300.000  5000.000 1410.000    61
+2.03599510E+01+2.36444020E-02-8.00996599E-06+1.23543694E-09-7.13457143E-14    2
-1.51264004E+04-7.57807484E+01+3.03844851E+00+6.35523371E-02-4.29455468E-05    3
+1.50665567E-08-2.16139351E-12-9.06691319E+03+1.74223348E+01+0.00000000E+00    4
C5H10O1-2  9/ 8/14      C   5H  10O   1    0G   300.000  5000.000 1424.000    31
+1.76453140E+01+2.17647043E-02-7.28831391E-06+1.11571673E-09-6.41056178E-14    2
-2.49627812E+04-6.94780751E+01-5.22384549E+00+7.95280569E-02-6.27918049E-05    3
+2.51187341E-08-3.99106436E-12-1.76152192E+04+5.15328120E+01+0.00000000E+00    4
C5H10O1-3  9/ 8/14      C   5H  10O   1    0G   300.000  5000.000 1445.000    21
+1.61536944E+01+2.22699220E-02-7.20967982E-06+1.07781327E-09-6.08828236E-14    2
-2.51216994E+04-6.18744318E+01-7.38770073E+00+8.62948016E-02-7.34565945E-05    3
+3.18221366E-08-5.43057938E-12-1.80648633E+04+6.09884425E+01+0.00000000E+00    4
C5H10O1-4  9/ 8/14      C   5H  10O   1    0G   300.000  5000.000 1470.000    11
+1.56838302E+01+2.28597182E-02-7.36869093E-06+1.09855828E-09-6.19425653E-14    2
-3.52365120E+04-6.06986511E+01-7.99511075E+00+8.48027993E-02-6.84820969E-05    3
+2.79646707E-08-4.48601572E-12-2.79347448E+04+6.36835324E+01+0.00000000E+00    4
C5H10O1-5  9/ 8/14      C   5H  10O   1    0G   300.000  5000.000 1447.000    01
+1.58722584E+01+2.41484940E-02-8.02830905E-06+1.22306406E-09-7.00384536E-14    2
-3.58667196E+04-6.73548909E+01-8.45066821E+00+8.36041573E-02-6.24375031E-05    3
+2.32498119E-08-3.38258239E-12-2.79060038E+04+6.19634163E+01+0.00000000E+00    4
C5H10O2-3  9/ 8/14      C   5H  10O   1    0G   300.000  5000.000 1415.000    31
+1.76695497E+01+2.16741351E-02-7.23760886E-06+1.10546424E-09-6.34044008E-14    2
-2.67999740E+04-7.01762004E+01-6.83688134E+00+9.00167224E-02-8.09486382E-05    3
+3.71523167E-08-6.73312332E-12-1.94907358E+04+5.73459463E+01+0.00000000E+00    4
C5H10O2-4  9/ 8/14      C   5H  10O   1    0G   300.000  5000.000 1396.000    21
+1.58873476E+01+2.48573824E-02-1.03962573E-05+1.95192708E-09-1.29464891E-13    2
-2.72224431E+04-6.26943208E+01-6.91381150E+00+8.65695113E-02-7.51445092E-05    3
+3.29307332E-08-5.77631101E-12-2.02336617E+04+5.66267224E+01+0.00000000E+00    4
C5H10OOH1-2O2 9/14      C   5H  11O   4    0G   300.000  5000.000 1394.000    71
+2.71105703E+01+2.34082367E-02-8.11719657E-06+1.27230537E-09-7.43221831E-14    2
-3.41406290E+04-1.08093476E+02+2.92123878E+00+7.67601721E-02-5.10111840E-05    3
+1.59643052E-08-1.82979631E-12-2.55486792E+04+2.27306226E+01+0.00000000E+00    4
C5H10OOH1-3O2 9/14      C   5H  11O   4    0G   300.000  5000.000 1394.000    71
+2.71105703E+01+2.34082367E-02-8.11719657E-06+1.27230537E-09-7.43221831E-14    2
-3.41406290E+04-1.08093476E+02+2.92123878E+00+7.67601721E-02-5.10111840E-05    3
+1.59643052E-08-1.82979631E-12-2.55486792E+04+2.27306226E+01+0.00000000E+00    4
C5H10OOH1-4O2 9/14      C   5H  11O   4    0G   300.000  5000.000 1394.000    71
+2.71105703E+01+2.34082367E-02-8.11719657E-06+1.27230537E-09-7.43221831E-14    2
-3.41406290E+04-1.08093476E+02+2.92123878E+00+7.67601721E-02-5.10111840E-05    3
+1.59643052E-08-1.82979631E-12-2.55486792E+04+2.27306226E+01+0.00000000E+00    4
C5H10OOH1-5O2 9/14      C   5H  11O   4    0G   300.000  5000.000 1390.000    71
+2.58212210E+01+2.46140917E-02-8.55565938E-06+1.34293065E-09-7.85178268E-14    2
-3.17158002E+04-9.97698267E+01+2.61115242E+00+7.58124541E-02-5.03939636E-05    3
+1.63241251E-08-2.04839461E-12-2.33970141E+04+2.58821117E+01+0.00000000E+00    4
C5H10OOH2-1O2 9/14      C   5H  11O   4    0G   300.000  5000.000 1394.000    71
+2.71105703E+01+2.34082367E-02-8.11719657E-06+1.27230537E-09-7.43221831E-14    2
-3.41406290E+04-1.08093476E+02+2.92123878E+00+7.67601721E-02-5.10111840E-05    3
+1.59643052E-08-1.82979631E-12-2.55486792E+04+2.27306226E+01+0.00000000E+00    4
C5H10OOH2-3O2 9/14      C   5H  11O   4    0G   300.000  5000.000 1405.000    71
+2.51554088E+01+2.42476887E-02-8.22109032E-06+1.26886123E-09-7.33157779E-14    2
-3.49522107E+04-9.69775586E+01+2.94958658E+00+7.94696642E-02-6.12300085E-05    3
+2.45360891E-08-3.99243941E-12-2.76263457E+04+2.10066180E+01+0.00000000E+00    4
C5H10OOH2-4O2 9/14      C   5H  11O   4    0G   300.000  5000.000 1405.000    71
+2.51554088E+01+2.42476887E-02-8.22109032E-06+1.26886123E-09-7.33157779E-14    2
-3.49522107E+04-9.69775586E+01+2.94958658E+00+7.94696642E-02-6.12300085E-05    3
+2.45360891E-08-3.99243941E-12-2.76263457E+04+2.10066180E+01+0.00000000E+00    4
C5H10OOH2-5O2 9/14      C   5H  11O   4    0G   300.000  5000.000 1394.000    71
+2.71105703E+01+2.34082367E-02-8.11719657E-06+1.27230537E-09-7.43221831E-14    2
-3.41406290E+04-1.08093476E+02+2.92123878E+00+7.67601721E-02-5.10111840E-05    3
+1.59643052E-08-1.82979631E-12-2.55486792E+04+2.27306226E+01+0.00000000E+00    4
C5H10OOH3-1O2 9/14      C   5H  11O   4    0G   300.000  5000.000 1394.000    71
+2.71105703E+01+2.34082367E-02-8.11719657E-06+1.27230537E-09-7.43221831E-14    2
-3.41406290E+04-1.08093476E+02+2.92123878E+00+7.67601721E-02-5.10111840E-05    3
+1.59643052E-08-1.82979631E-12-2.55486792E+04+2.27306226E+01+0.00000000E+00    4
C5H10OOH3-2O2 9/14      C   5H  11O   4    0G   300.000  5000.000 1405.000    71
+2.51554088E+01+2.42476887E-02-8.22109032E-06+1.26886123E-09-7.33157779E-14    2
-3.49522107E+04-9.69775586E+01+2.94958658E+00+7.94696642E-02-6.12300085E-05    3
+2.45360891E-08-3.99243941E-12-2.76263457E+04+2.10066180E+01+0.00000000E+00    4
C5H91-2,3OOH  9/14      C   5H  11O   4    0G   300.000  5000.000 1405.000    81
+2.55056147E+01+2.36990320E-02-8.07032909E-06+1.24934920E-09-7.23427367E-14    2
-2.71353489E+04-9.69348818E+01+2.91226160E+00+7.95651114E-02-6.13230261E-05    3
+2.44460527E-08-3.95034020E-12-1.96516956E+04+2.32188202E+01+0.00000000E+00    4
C5H91-2,4OOH  9/14      C   5H  11O   4    0G   300.000  5000.000 1405.000    81
+2.55056147E+01+2.36990320E-02-8.07032909E-06+1.24934920E-09-7.23427367E-14    2
-2.71353489E+04-9.69348818E+01+2.91226160E+00+7.95651114E-02-6.13230261E-05    3
+2.44460527E-08-3.95034020E-12-1.96516956E+04+2.32188202E+01+0.00000000E+00    4
C5H91-2,5OOH  9/14      C   5H  11O   4    0G   300.000  5000.000 1397.000    81
+2.50741397E+01+2.44380043E-02-8.40704928E-06+1.31038422E-09-7.62381905E-14    2
-2.51871158E+04-9.38667514E+01+2.56086129E+00+7.80408775E-02-5.74863330E-05    3
+2.18761227E-08-3.39924240E-12-1.74851061E+04+2.66588551E+01+0.00000000E+00    4
C5H91-3,4OOH  9/14      C   5H  11O   4    0G   300.000  5000.000 1405.000    81
+2.54680852E+01+2.36307420E-02-8.02474436E-06+1.23994908E-09-7.17032304E-14    2
-2.70635665E+04-9.67605580E+01+2.48775154E+00+8.15271831E-02-6.44013124E-05    3
+2.63443736E-08-4.35804025E-12-1.95635349E+04+2.50626503E+01+0.00000000E+00    4
C5H91-3,5OOH  9/14      C   5H  11O   4    0G   300.000  5000.000 1397.000    81
+2.75716451E+01+2.26282394E-02-7.85651555E-06+1.23251566E-09-7.20426920E-14    2
-2.62702922E+04-1.08648340E+02+2.50132978E+00+7.93141150E-02-5.51608762E-05    3
+1.83963651E-08-2.32880956E-12-1.75129588E+04+2.64329747E+01+0.00000000E+00    4
C5H91-4,5OOH  9/14      C   5H  11O   4    0G   300.000  5000.000 1397.000    81
+2.75716451E+01+2.26282394E-02-7.85651555E-06+1.23251566E-09-7.20426920E-14    2
-2.62702922E+04-1.08648340E+02+2.50132978E+00+7.93141150E-02-5.51608762E-05    3
+1.83963651E-08-2.32880956E-12-1.75129588E+04+2.64329747E+01+0.00000000E+00    4
C5H92-1,3OOH  9/14      C   5H  11O   4    0G   300.000  5000.000 1413.000    81
+2.46778451E+01+2.47896676E-02-8.53168232E-06+1.33018418E-09-7.74050315E-14    2
-2.64008851E+04-9.18794025E+01+3.42922915E+00+7.33174178E-02-5.05533009E-05    3
+1.77709491E-08-2.53421378E-12-1.89212844E+04+2.26144479E+01+0.00000000E+00    4
C5H92-1,4OOH  9/14      C   5H  11O   4    0G   300.000  5000.000 1413.000    81
+2.46778451E+01+2.47896676E-02-8.53168232E-06+1.33018418E-09-7.74050315E-14    2
-2.64008851E+04-9.18794025E+01+3.42922915E+00+7.33174178E-02-5.05533009E-05    3
+1.77709491E-08-2.53421378E-12-1.89212844E+04+2.26144479E+01+0.00000000E+00    4
C5H92-1,5OOH  9/14      C   5H  11O   4    0G   300.000  5000.000 1399.000    81
+2.63836136E+01+2.38373273E-02-8.31679219E-06+1.30877666E-09-7.66591074E-14    2
-2.52930801E+04-1.01118754E+02+3.43107332E+00+7.25133538E-02-4.53395240E-05    3
+1.29499313E-08-1.26534785E-12-1.69000809E+04+2.37843821E+01+0.00000000E+00    4
C5H92-3,4OOH  9/14      C   5H  11O   4    0G   300.000  5000.000 1418.000    81
+2.51070211E+01+2.40686276E-02-8.20467040E-06+1.27103065E-09-7.36339262E-14    2
-2.83591157E+04-9.49637963E+01+3.76788328E+00+7.47668469E-02-5.41780015E-05    3
+2.01841133E-08-3.04867679E-12-2.10823293E+04+1.92561961E+01+0.00000000E+00    4
C5H92-3,5OOH  9/14      C   5H  11O   4    0G   300.000  5000.000 1413.000    81
+2.46778451E+01+2.47896676E-02-8.53168232E-06+1.33018418E-09-7.74050315E-14    2
-2.64008851E+04-9.18794025E+01+3.42922915E+00+7.33174178E-02-5.05533009E-05    3
+1.77709491E-08-2.53421378E-12-1.89212844E+04+2.26144479E+01+0.00000000E+00    4
C5H92-4,5OOH  9/14      C   5H  11O   4    0G   300.000  5000.000 1413.000    81
+2.47514622E+01+2.41459993E-02-8.18238994E-06+1.26250806E-09-7.29352454E-14    2
-2.63782993E+04-9.11444444E+01+4.06621416E+00+7.20273834E-02-4.95956461E-05    3
+1.70908613E-08-2.31584179E-12-1.92523266E+04+1.99316930E+01+0.00000000E+00    4
C5H93-1,2OOH  9/14      C   5H  11O   4    0G   300.000  5000.000 1413.000    81
+2.46778451E+01+2.47896676E-02-8.53168232E-06+1.33018418E-09-7.74050315E-14    2
-2.64008851E+04-9.18794025E+01+3.42922915E+00+7.33174178E-02-5.05533009E-05    3
+1.77709491E-08-2.53421378E-12-1.89212844E+04+2.26144479E+01+0.00000000E+00    4
C5H93-1,4OOH  9/14      C   5H  11O   4    0G   300.000  5000.000 1413.000    81
+2.46778451E+01+2.47896676E-02-8.53168232E-06+1.33018418E-09-7.74050315E-14    2
-2.64008851E+04-9.18794025E+01+3.42922915E+00+7.33174178E-02-5.05533009E-05    3
+1.77709491E-08-2.53421378E-12-1.89212844E+04+2.26144479E+01+0.00000000E+00    4
C5H93-1,5OOH  9/14      C   5H  11O   4    0G   300.000  5000.000 1399.000    81
+2.44184921E+01+2.49501505E-02-8.57440942E-06+1.33558596E-09-7.76697869E-14    2
-2.45529807E+04-8.95288488E+01+3.67511835E+00+6.98557277E-02-4.39193701E-05    3
+1.31290152E-08-1.43358803E-12-1.70587842E+04+2.30262907E+01+0.00000000E+00    4
C5H93-2,4OOH  9/14      C   5H  11O   4    0G   300.000  5000.000 1418.000    81
+2.51070211E+01+2.40686276E-02-8.20467040E-06+1.27103065E-09-7.36339262E-14    2
-2.83591157E+04-9.56532779E+01+3.76788328E+00+7.47668469E-02-5.41780015E-05    3
+2.01841133E-08-3.04867679E-12-2.10823293E+04+1.85667144E+01+0.00000000E+00    4
C5H91-3OOH  9/8/14      C   5H  10O   2    0G   300.000  5000.000 1394.000    51
+2.24660467E+01+2.00408413E-02-6.84550040E-06+1.06266050E-09-6.16741604E-14    2
-2.26148518E+04-9.04469895E+01-1.89589507E+00+8.18483531E-02-6.75161021E-05    3
+2.83331852E-08-4.76826956E-12-1.47140793E+04+3.85399143E+01+0.00000000E+00    4
C5H91-4OOH  9/8/14      C   5H  10O   2    0G   300.000  5000.000 1402.000    51
+1.96307052E+01+2.22000091E-02-7.52489271E-06+1.16109117E-09-6.70722374E-14    2
-2.30400033E+04-7.32135194E+01+1.38243484E+00+6.67661361E-02-4.96344237E-05    3
+1.94278468E-08-3.12175781E-12-1.69086691E+04+2.40815942E+01+0.00000000E+00    4
C5H91-5OOH  9/8/14      C   5H  10O   2    0G   300.000  5000.000 1392.000    51
+1.93103284E+01+2.29913370E-02-7.91269843E-06+1.23358507E-09-7.17773402E-14    2
-2.12246688E+04-7.09825558E+01+9.93373748E-01+6.46025217E-02-4.40191862E-05    3
+1.55375290E-08-2.26236370E-12-1.47156820E+04+2.78588419E+01+0.00000000E+00    4
C5H92-1OOH  9/8/14      C   5H  10O   2    0G   300.000  5000.000 1382.000    51
+2.10623695E+01+2.15772208E-02-7.44876502E-06+1.16423903E-09-6.78819533E-14    2
-2.15816942E+04-8.04705541E+01+5.77880009E-01+6.91528527E-02-5.00924279E-05    3
+1.88100079E-08-2.91765412E-12-1.44043272E+04+2.97056559E+01+0.00000000E+00    4
C5H92-4OOH  9/8/14      C   5H  10O   2    0G   300.000  5000.000 1389.000    51
+2.22714879E+01+1.99891269E-02-6.78760139E-06+1.05004677E-09-6.08129638E-14    2
-2.39098291E+04-9.00213678E+01-1.10664142E+00+7.70652343E-02-6.01781689E-05    3
+2.37846489E-08-3.77298555E-12-1.61217479E+04+3.45219377E+01+0.00000000E+00    4
C5H92-5OOH  9/8/14      C   5H  10O   2    0G   300.000  5000.000 1389.000    51
+1.88657282E+01+2.33222202E-02-8.01683595E-06+1.24882522E-09-7.26244846E-14    2
-2.24129903E+04-6.91316665E+01+1.76944896E+00+6.00153444E-02-3.72031347E-05    3
+1.14551487E-08-1.39226390E-12-1.61243818E+04+2.38818885E+01+0.00000000E+00    4
C5H9O1-2OOH-3 9/14      C   5H  10O   3    0G   300.000  5000.000 1422.000    51
+2.40742385E+01+2.10049879E-02-7.12965508E-06+1.10196053E-09-6.37577378E-14    2
-3.86905727E+04-9.86614868E+01-1.63458528E+00+8.37428576E-02-6.46448858E-05    3
+2.45435115E-08-3.63637746E-12-3.02443795E+04+3.81009801E+01+0.00000000E+00    4
C5H9O1-2OOH-4 9/14      C   5H  10O   3    0G   300.000  5000.000 1422.000    51
+2.40742385E+01+2.10049879E-02-7.12965508E-06+1.10196053E-09-6.37577378E-14    2
-3.86905727E+04-9.86614868E+01-1.63458528E+00+8.37428576E-02-6.46448858E-05    3
+2.45435115E-08-3.63637746E-12-3.02443795E+04+3.81009801E+01+0.00000000E+00    4
C5H9O1-2OOH-5 9/14      C   5H  10O   3    0G   300.000  5000.000 1425.000    51
+2.31521586E+01+2.15716913E-02-7.27787584E-06+1.12021946E-09-6.46248595E-14    2
-3.63754336E+04-9.23672941E+01-2.91502569E+00+8.63720024E-02-6.80858869E-05    3
+2.66150873E-08-4.08265327E-12-2.79298051E+04+4.58804153E+01+0.00000000E+00    4
C5H9O1-3OOH-2 9/14      C   5H  10O   3    0G   300.000  5000.000 1421.000    41
+2.29238871E+01+2.22244781E-02-7.50929996E-06+1.15689292E-09-6.67794310E-14    2
-3.93149495E+04-9.38426660E+01-4.67708778E+00+9.25191737E-02-7.56245586E-05    3
+3.08655754E-08-4.96974700E-12-3.05178886E+04+5.19807893E+01+0.00000000E+00    4
C5H9O1-3OOH-4 9/14      C   5H  10O   3    0G   300.000  5000.000 1421.000    41
+2.29238871E+01+2.22244781E-02-7.50929996E-06+1.15689292E-09-6.67794310E-14    2
-3.93149495E+04-9.38426660E+01-4.67708778E+00+9.25191737E-02-7.56245586E-05    3
+3.08655754E-08-4.96974700E-12-3.05178886E+04+5.19807893E+01+0.00000000E+00    4
C5H9O1-3OOH-5 9/14      C   5H  10O   3    0G   300.000  5000.000 1421.000    41
+2.21702811E+01+2.28760461E-02-7.73630997E-06+1.19254044E-09-6.88630410E-14    2
-3.71502930E+04-8.87113724E+01-5.55071358E+00+9.29081113E-02-7.49705054E-05    3
+3.02210571E-08-4.80852681E-12-2.82561346E+04+5.79510604E+01+0.00000000E+00    4
C5H9O1-4OOH-2 9/14      C   5H  10O   3    0G   300.000  5000.000 1417.000    31
+2.17260410E+01+2.34146274E-02-7.86187868E-06+1.20571561E-09-6.93653621E-14    2
-4.90509096E+04-8.83590566E+01-9.18084516E+00+1.08786371E-01-9.86756121E-05    3
+4.49207522E-08-8.03087742E-12-3.98013189E+04+7.26760969E+01+0.00000000E+00    4
C5H9O1-4OOH-3 9/14      C   5H  10O   3    0G   300.000  5000.000 1417.000    31
+2.17260410E+01+2.34146274E-02-7.86187868E-06+1.20571561E-09-6.93653621E-14    2
-4.90509096E+04-8.83590566E+01-9.18084516E+00+1.08786371E-01-9.86756121E-05    3
+4.49207522E-08-8.03087742E-12-3.98013189E+04+7.26760969E+01+0.00000000E+00    4
C5H9O1-4OOH-5 9/14      C   5H  10O   3    0G   300.000  5000.000 1411.000    31
+2.13868464E+01+2.42467386E-02-8.26745278E-06+1.28123479E-09-7.42527951E-14    2
-4.72411464E+04-8.60552096E+01-9.29661331E+00+1.04958911E-01-9.00892767E-05    3
+3.89843596E-08-6.68819849E-12-3.76382956E+04+7.52773731E+01+0.00000000E+00    4
C5H9O1-5OOH-2 9/14      C   5H  10O   3    0G   300.000  5000.000 1407.000    21
+2.24618796E+01+2.42252273E-02-8.36381388E-06+1.30712783E-09-7.62010208E-14    2
-5.00102121E+04-9.76835754E+01-9.63082131E+00+1.06539535E-01-8.95953916E-05    3
+3.77712411E-08-6.32248900E-12-3.97499469E+04+7.18166046E+01+0.00000000E+00    4
C5H9O1-5OOH-3 9/14      C   5H  10O   3    0G   300.000  5000.000 1407.000    21
+2.24618796E+01+2.42252273E-02-8.36381388E-06+1.30712783E-09-7.62010208E-14    2
-5.00102121E+04-9.83780898E+01-9.63082131E+00+1.06539535E-01-8.95953916E-05    3
+3.77712411E-08-6.32248900E-12-3.97499469E+04+7.11220903E+01+0.00000000E+00    4
C5H9O2-3OOH-1 9/14      C   5H  10O   3    0G   300.000  5000.000 1436.000    51
+2.37309690E+01+2.06751517E-02-6.88444402E-06+1.05044759E-09-6.02362275E-14    2
-3.84362991E+04-9.61945548E+01-2.95211763E+00+8.90845071E-02-7.32339295E-05    3
+2.98425405E-08-4.76173344E-12-3.00280666E+04+4.45334764E+01+0.00000000E+00    4
C5H9O2-3OOH-4 9/14      C   5H  10O   3    0G   300.000  5000.000 1430.000    51
+2.36691815E+01+1.92560232E-02-6.07856844E-06+8.92371727E-10-4.97448691E-14    2
-3.96296162E+04-9.51544015E+01-4.57026018E+00+1.05196229E-01-1.05063534E-04    3
+5.15547206E-08-9.70822253E-12-3.20442434E+04+4.90445735E+01+0.00000000E+00    4
C5H9O2-3OOH-5 9/14      C   5H  10O   3    0G   300.000  5000.000 1436.000    51
+2.37309690E+01+2.06751517E-02-6.88444402E-06+1.05044759E-09-6.02362275E-14    2
-3.84362991E+04-9.61945548E+01-2.95211763E+00+8.90845071E-02-7.32339295E-05    3
+2.98425405E-08-4.76173344E-12-3.00280666E+04+4.45334764E+01+0.00000000E+00    4
C5H9O2-4OOH-1 9/14      C   5H  10O   3    0G   300.000  5000.000 1429.000    41
+2.26534501E+01+2.20609304E-02-7.36975144E-06+1.12674313E-09-6.46941132E-14    2
-3.91616134E+04-9.19653554E+01-5.54951868E+00+9.55182117E-02-8.01619637E-05    3
+3.35588175E-08-5.52327105E-12-3.03610773E+04+5.64175360E+01+0.00000000E+00    4
C5H9O2-4OOH-3 9/14      C   5H  10O   3    0G   300.000  5000.000 1427.000    41
+2.36121225E+01+2.13802117E-02-7.16433060E-06+1.09773009E-09-6.31280098E-14    2
-4.14634634E+04-9.91050535E+01-4.69459258E+00+9.49457030E-02-7.98763001E-05    3
+3.34048886E-08-5.48568419E-12-3.26159152E+04+4.98789194E+01+0.00000000E+00    4
C5H9O1-2O-5 9/8/14      C   5H   9O   2    0G   300.000  5000.000 1421.000    31
+2.01220485E+01+2.03728898E-02-6.96642194E-06+1.08201705E-09-6.28152071E-14    2
-1.74886279E+04-7.89086914E+01-6.46243908E-01+6.53341554E-02-4.13295267E-05    3
+1.15534981E-08-9.90013428E-13-1.01037208E+04+3.35841975E+01+0.00000000E+00    4
CH2CH2OCH2CH2CHO 4      C   5H   9O   2    0G   300.000  5000.000 1447.000    51
+1.75698412E+01+2.05459822E-02-6.77593971E-06+1.02644892E-09-5.85405221E-14    2
-2.62366696E+04-5.93672925E+01-6.18508829E-01+6.43128028E-02-4.60370456E-05    3
+1.65228932E-08-2.31382679E-12-2.02103439E+04+3.75876155E+01+0.00000000E+00    4
NC5KET12   9/ 8/14      C   5H  10O   3    0G   300.000  5000.000 1386.000    61
+2.56958620E+01+1.97581564E-02-6.83008913E-06+1.06937987E-09-6.24522080E-14    2
-4.91027960E+04-1.03505108E+02-1.29174799E+00+8.64138926E-02-7.02456071E-05    3
+2.86657248E-08-4.68321816E-12-4.01718501E+04+4.00248297E+01+0.00000000E+00    4
NC5KET13   9/ 8/14      C   5H  10O   3    0G   300.000  5000.000 1405.000    61
+2.25901874E+01+2.17812117E-02-7.38063794E-06+1.13910638E-09-6.58295642E-14    2
-4.92679139E+04-8.65971472E+01+3.00527399E+00+6.57859047E-02-4.36348536E-05    3
+1.39803001E-08-1.68002311E-12-4.24094861E+04+1.90078452E+01+0.00000000E+00    4
NC5KET14   9/ 8/14      C   5H  10O   3    0G   300.000  5000.000 1405.000    61
+2.25901874E+01+2.17812117E-02-7.38063794E-06+1.13910638E-09-6.58295642E-14    2
-4.92679139E+04-8.65971472E+01+3.00527399E+00+6.57859047E-02-4.36348536E-05    3
+1.39803001E-08-1.68002311E-12-4.24094861E+04+1.90078452E+01+0.00000000E+00    4
NC5KET15   9/ 8/14      C   5H  10O   3    0G   300.000  5000.000 1389.000    61
+2.22256536E+01+2.26347088E-02-7.79347724E-06+1.21574025E-09-7.07808477E-14    2
-4.74266046E+04-8.41025053E+01+2.63079123E+00+6.36042087E-02-3.80050385E-05    3
+1.00772174E-08-8.15255520E-13-4.02201480E+04+2.27068767E+01+0.00000000E+00    4
NC5KET21   9/ 8/14      C   5H  10O   3    0G   300.000  5000.000 1388.000    61
+2.45822715E+01+2.02064434E-02-6.87782149E-06+1.06593008E-09-6.18171916E-14    2
-5.02288346E+04-9.64925259E+01-1.97528990E-01+7.92952922E-02-6.01376298E-05    3
+2.26192730E-08-3.36572580E-12-4.18751690E+04+3.59471835E+01+0.00000000E+00    4
NC5KET23   9/ 8/14      C   5H  10O   3    0G   300.000  5000.000 1390.000    61
+2.42608382E+01+2.03281864E-02-6.88576173E-06+1.06357099E-09-6.15324796E-14    2
-5.21063936E+04-9.49416999E+01-4.59062579E-01+8.23364070E-02-6.69200221E-05    3
+2.76548457E-08-4.58692734E-12-4.40257491E+04+3.61810105E+01+0.00000000E+00    4
NC5KET24   9/ 8/14      C   5H  10O   3    0G   300.000  5000.000 1417.000    61
+2.13557506E+01+2.20059280E-02-7.28286282E-06+1.10610540E-09-6.32057101E-14    2
-5.23446138E+04-7.91468873E+01+3.70377687E+00+6.22140345E-02-4.08903819E-05    3
+1.31907442E-08-1.60742182E-12-4.62411438E+04+1.58017148E+01+0.00000000E+00    4
NC5KET25   9/ 8/14      C   5H  10O   3    0G   300.000  5000.000 1395.000    61
+2.09051806E+01+2.29956432E-02-7.75343394E-06+1.19262969E-09-6.87612656E-14    2
-5.04678003E+04-7.61623703E+01+3.30376112E+00+6.01763378E-02-3.55337358E-05    3
+9.49960340E-09-7.96339342E-13-4.40485734E+04+1.96186974E+01+0.00000000E+00    4
NC5KET31   9/ 8/14      C   5H  10O   3    0G   300.000  5000.000 1431.000    61
+2.14962676E+01+2.20658980E-02-7.35490387E-06+1.12358588E-09-6.45028163E-14    2
-5.08471346E+04-8.02429953E+01+4.06393861E+00+5.46274576E-02-2.50666165E-05    3
+2.02312915E-09+1.00150274E-12-4.41625000E+04+1.59654525E+01+0.00000000E+00    4
NC5KET32   9/ 8/14      C   5H  10O   3    0G   300.000  5000.000 1388.000    61
+2.43326367E+01+2.02926765E-02-6.88030752E-06+1.06352004E-09-6.15648338E-14    2
-5.22889844E+04-9.61325613E+01+3.80342038E-01+7.67072849E-02-5.67635185E-05    3
+2.07068449E-08-2.96497951E-12-4.41579478E+04+3.21097700E+01+0.00000000E+00    4
NC5KET12O  9/ 8/14      C   5H   9O   2    0G   300.000  5000.000 1377.000    41
+2.09367959E+01+2.00874425E-02-7.04829670E-06+1.11330293E-09-6.53771464E-14    2
-3.04314417E+04-8.04081881E+01+2.82328315E+00+5.56013887E-02-3.02956498E-05    3
+6.22735484E-09-8.25379616E-14-2.35055878E+04+1.92120018E+01+0.00000000E+00    4
NC5KET13O  9/ 8/14      C   5H   9O   2    0G   300.000  5000.000 1323.000    41
+2.11225120E+01+1.90830240E-02-6.52403075E-06+1.01368310E-09-5.88793478E-14    2
-3.11151636E+04-8.21812017E+01+3.92095399E+00+4.94038774E-02-1.99599619E-05    3
-1.05666833E-09+1.70331197E-12-2.43649054E+04+1.33502699E+01+0.00000000E+00    4
NC5KET14O  9/ 8/14      C   5H   9O   2    0G   300.000  5000.000 1323.000    41
+2.11225120E+01+1.90830240E-02-6.52403075E-06+1.01368310E-09-5.88793478E-14    2
-3.11151636E+04-8.21812017E+01+3.92095399E+00+4.94038774E-02-1.99599619E-05    3
-1.05666833E-09+1.70331197E-12-2.43649054E+04+1.33502699E+01+0.00000000E+00    4
NC5KET15O  9/ 8/14      C   5H   9O   2    0G   300.000  5000.000 1489.000    41
+1.92273388E+01+2.11348590E-02-7.32088660E-06+1.14667396E-09-6.69507752E-14    2
-2.85866827E+04-7.08964819E+01+3.41522476E+00+4.72023685E-02-1.66453220E-05    3
-2.39548810E-09+1.83814508E-12-2.21147912E+04+1.77035103E+01+0.00000000E+00    4
NC5KET21O  9/ 8/14      C   5H   9O   2    0G   300.000  5000.000 1669.000    41
+1.55374345E+01+2.65967153E-02-9.82520086E-06+1.61087197E-09-9.71864472E-14    2
-2.96220202E+04-4.97983106E+01+7.57725086E+00+3.09672386E-02+2.94905694E-06    3
-1.10969895E-08+3.01674992E-12-2.56340563E+04-2.16720088E+00+0.00000000E+00    4
NC5KET23O  9/ 8/14      C   5H   9O   2    0G   300.000  5000.000 1383.000    41
+1.95245872E+01+2.08858647E-02-7.23257140E-06+1.13238277E-09-6.60902126E-14    2
-3.34926354E+04-7.21145428E+01+3.56460361E+00+5.18213432E-02-2.70330790E-05    3
+5.19426451E-09+1.69499746E-14-2.73448675E+04+1.58030522E+01+0.00000000E+00    4
NC5KET24O  9/ 8/14      C   5H   9O   2    0G   300.000  5000.000 1382.000    41
+1.87900628E+01+2.10010240E-02-7.16188369E-06+1.11001257E-09-6.43339326E-14    2
-3.32898658E+04-6.78862933E+01+4.40946289E+00+4.75586902E-02-2.19238261E-05    3
+2.43250490E-09+5.88504938E-13-2.76535939E+04+1.17394140E+01+0.00000000E+00    4
NC5KET25O  9/ 8/14      C   5H   9O   2    0G   300.000  5000.000 1433.000    41
+1.81303967E+01+2.13611121E-02-7.24506108E-06+1.11897303E-09-6.47006005E-14    2
-3.16682816E+04-6.41505194E+01+4.40785464E+00+4.34772079E-02-1.40284695E-05    3
-3.02310104E-09+1.86768676E-12-2.60265017E+04+1.28766258E+01+0.00000000E+00    4
NC5KET31O  9/ 8/14      C   5H   9O   2    0G   300.000  5000.000 1426.000    41
+1.92416140E+01+2.07624762E-02-7.12773261E-06+1.11092657E-09-6.46775655E-14    2
-3.25710561E+04-7.19638232E+01+5.37524822E+00+3.49659305E-02+3.67920037E-06    3
-1.56750631E-08+4.84743343E-12-2.61248405E+04+8.64755527E+00+0.00000000E+00    4
NC5KET32O  9/ 8/14      C   5H   9O   2    0G   300.000  5000.000 1539.000    41
+1.90206162E+01+2.10022758E-02-7.20628551E-06+1.12155484E-09-6.51936687E-14    2
-3.33553472E+04-6.97524186E+01+4.55782533E+00+4.55546283E-02-1.73485031E-05    3
-9.24152417E-10+1.38889438E-12-2.74919397E+04+1.10596626E+01+0.00000000E+00    4
NC5DIONE13  10/15  THERMC   5H   8O   2    0G   300.000  5000.000 1380.000    41
+1.81672199E+01+1.95477748E-02-6.78556722E-06+1.06428037E-09-6.21973311E-14    2
-5.11134997E+04-6.80388452E+01+1.16337913E+00+5.32067868E-02-2.90297512E-05    3
+5.99807535E-09-7.60467747E-14-4.46714058E+04+2.53180917E+01+0.00000000E+00    4
NC5DIONE24  10/15  THERMC   5H   8O   2    0G   300.000  5000.000 1393.000    41
+1.63259547E+01+2.07678096E-02-7.12494176E-06+1.10833798E-09-6.43882952E-14    2
-5.38361320E+04-5.71667682E+01+1.23573850E+00+5.44884679E-02-3.57895292E-05    3
+1.21944125E-08-1.71810392E-12-4.84057706E+04+2.44807388E+01+0.00000000E+00    4
C5H10OH23  9/ 8/14      C   5H  11O   1    0G   300.000  5000.000 1447.000    51
+1.70150141E+01+2.35005444E-02-7.77847758E-06+1.18102788E-09-6.74584591E-14    2
-2.30013982E+04-5.87178603E+01+9.23102001E-01+5.84732430E-02-3.47946675E-05    3
+9.61256846E-09-8.64039220E-13-1.72758426E+04+2.84227761E+01+0.00000000E+00    4
O2C5H10OH23 9/8/14      C   5H  11O   3    0G   300.000  5000.000 1413.000    61
+2.25663309E+01+2.36960784E-02-7.89320309E-06+1.20343029E-09-6.89316529E-14    2
-4.25964462E+04-8.48729630E+01+1.48292990E+00+7.92100619E-02-6.45238925E-05    3
+2.75597603E-08-4.74651399E-12-3.59663215E+04+2.60236189E+01+0.00000000E+00    4
OCH2CHO    9/ 8/14      C   2H   3O   2    0G   300.000  5000.000 1468.000    11
+9.83472746E+00+7.77895515E-03-2.78174926E-06+4.44911597E-10-2.63530280E-14    2
-1.50740413E+04-2.41644767E+01+6.12784775E+00+6.67998271E-03+1.00125301E-05    3
-1.06887671E-08+2.76652784E-12-1.28216539E+04-8.09763223E-01+0.00000000E+00    4
CH2OCH2CHO 9/ 8/14      C   3H   5O   2    0G   300.000  5000.000 1386.000    31
+1.11192754E+01+1.27912900E-02-4.35464414E-06+6.73922275E-10-3.90118722E-14    2
-1.79694096E+04-2.74688068E+01+4.09796526E+00+2.50971166E-02-1.04380487E-05    3
+6.95156168E-10+3.93228907E-13-1.51203149E+04+1.16942054E+01+0.00000000E+00    4
C2H4OCHO   9/ 8/14      C   3H   5O   2    0G   300.000  5000.000 1684.000    21
+1.22682078E+01+1.37336751E-02-5.06732537E-06+8.30265992E-10-5.00728023E-14    2
-2.09125606E+04-3.56985038E+01+3.11985293E+00+3.19514120E-02-1.67508873E-05    3
+3.25914973E-09-4.96818754E-14-1.76239471E+04+1.42845094E+01+0.00000000E+00    4
C5H10OOH1-3OH  10/14/15 C   5H  12O   3    0G   300.000  5000.000 1403.000    71
+2.31192753E+01+2.59986683E-02-8.82860426E-06+1.36395720E-09-7.88606733E-14    2
-5.79892376E+04-8.81999105E+01+3.54670341E-01+8.27825400E-02-6.38327513E-05    3
+2.58589986E-08-4.28053334E-12-5.04620388E+04+3.27492018E+01+0.00000000E+00    4
C5H10OOH2-4OH  10/14/15 C   5H  12O   3    0G   300.000  5000.000 1411.000    71
+2.35162773E+01+2.51435990E-02-8.42079438E-06+1.28867610E-09-7.40107760E-14    2
-5.98557610E+04-9.09142876E+01+7.69420941E-01+8.47002755E-02-6.89331076E-05    3
+2.93938563E-08-5.06044347E-12-5.26556407E+04+2.88739602E+01+0.00000000E+00    4
C5H10OOH3-1OH  10/14/15 C   5H  12O   3    0G   300.000  5000.000 1406.000    71
+2.38716811E+01+2.53396515E-02-8.59895412E-06+1.32803347E-09-7.67709894E-14    2
-5.82703781E+04-9.26845624E+01+7.53538721E-01+8.16716738E-02-6.11918401E-05    3
+2.36490302E-08-3.69940856E-12-5.05457936E+04+3.05276339E+01+0.00000000E+00    4
NC5CYCPER13  11/15 THERMC   5H  10O   3    0G   300.000  5000.000 1407.000    31
+2.41561308E+01+2.24095731E-02-7.74873939E-06+1.21233645E-09-7.07323367E-14    2
-5.55344567E+04-1.03522127E+02-4.99453890E+00+9.45988114E-02-7.58465481E-05    3
+3.02152876E-08-4.76416624E-12-4.59881161E+04+5.13024248E+01+0.00000000E+00    4
NC5CYCPER24  11/15 THERMC   5H  10O   3    0G   300.000  5000.000 1408.000    31
+2.22820691E+01+2.33310062E-02-7.91636135E-06+1.22269476E-09-7.06906786E-14    2
-5.60698326E+04-9.35418515E+01-4.25869873E+00+9.26924392E-02-7.79864322E-05    3
+3.34971276E-08-5.74390775E-12-4.76901635E+04+4.62163973E+01+0.00000000E+00    4
NC5CYCPER31  11/15 THERMC   5H  10O   3    0G   300.000  5000.000 1400.000    31
+2.20861156E+01+2.39837041E-02-8.24798762E-06+1.28546679E-09-7.47886437E-14    2
-5.42162418E+04-9.20233359E+01-4.01647605E+00+8.90855731E-02-7.09557408E-05    3
+2.89246712E-08-4.75384108E-12-4.56274320E+04+4.65938612E+01+0.00000000E+00    4
IC5H12     17/8/15      C   5H  12    0    0G   300.000  5000.000 1397.000    41
+1.58024165E+01+2.58962455E-02-8.80211277E-06+1.36051024E-09-7.86804753E-14    2
-2.64876700E+04-6.08691324E+01-1.61700908E+00+6.68962508E-02-4.65394790E-05    3
+1.75637406E-08-2.80513304E-12-2.03922408E+04+3.27016966E+01+0.00000000E+00    4
AC5H11     17/8/15      C   5H  11    0    0G   300.000  5000.000 1397.000    41
+1.52292407E+01+2.38482717E-02-8.09849455E-06+1.25096662E-09-7.23133933E-14    2
-1.35828406E+03-5.42832371E+01-1.22777654E+00+6.32926027E-02-4.52076107E-05    3
+1.75515079E-08-2.87257258E-12+4.32562497E+03+3.38598206E+01+0.00000000E+00    4
BC5H11     17/8/15      C   5H  11    0    0G   300.000  5000.000 1385.000    41
+1.41464948E+01+2.48340049E-02-8.45503425E-06+1.30848803E-09-7.57429130E-14    2
-3.88001657E+03-4.87192778E+01+1.65843160E+00+4.60868150E-02-1.82956944E-05    3
+8.82319315E-10+7.56537666E-13+1.29054584E+03+2.12275239E+01+0.00000000E+00    4
CC5H11     17/8/15      C   5H  11    0    0G   300.000  5000.000 1402.000    41
+1.43628831E+01+2.43459715E-02-8.21904266E-06+1.26457869E-09-7.28991288E-14    2
-2.64593539E+03-4.96386458E+01+1.97886349E-01+5.35219440E-02-2.95961594E-05    3
+7.61177489E-09-6.45328560E-13+2.66542853E+03+2.78232188E+01+0.00000000E+00    4
DC5H11     17/8/15      C   5H  11    0    0G   300.000  5000.000 1397.000    41
+1.52292407E+01+2.38482717E-02-8.09849455E-06+1.25096662E-09-7.23133933E-14    2
-1.35828406E+03-5.49727188E+01-1.22777654E+00+6.32926027E-02-4.52076107E-05    3
+1.75515079E-08-2.87257258E-12+4.32562497E+03+3.31703389E+01+0.00000000E+00    4
AC5H9O-A2  9/ 8/14      C   5H   9O   1    0G   300.000  5000.000 1364.000    31
+1.67516787E+01+2.16463662E-02-7.61269705E-06+1.20404408E-09-7.07632803E-14    2
-3.95848360E+03-6.08201916E+01+4.66263417E+00+3.89775126E-02-1.12815501E-05    3
-2.66550677E-09+1.40115432E-12+1.47086581E+03+8.21346271E+00+0.00000000E+00    4
AC5H11O2H  17/8/15      C   5H  12O   2    0G   300.000  5000.000 1397.000    61
+2.08513274E+01+2.60811030E-02-8.91735578E-06+1.38397232E-09-8.02716539E-14    2
-3.77194279E+04-8.04522304E+01-4.76374815E-01+7.83789321E-02-5.91712555E-05    3
+2.38263919E-08-3.97732270E-12-3.05087904E+04+3.32977557E+01+0.00000000E+00    4
BC5H11O2H  17/8/15      C   5H  12O   2    0G   300.000  5000.000 1389.000    61
+2.07291068E+01+2.60358698E-02-8.86783077E-06+1.37263265E-09-7.94629195E-14    2
-4.16991829E+04-8.29348605E+01+7.48347855E-01+7.54437451E-02-5.69961198E-05    3
+2.32342064E-08-3.94363492E-12-3.49638594E+04+2.35201019E+01+0.00000000E+00    4
CC5H11O2H  17/8/15      C   5H  12O   2    0G   300.000  5000.000 1406.000    61
+2.11504126E+01+2.53098885E-02-8.53703900E-06+1.31271216E-09-7.56412244E-14    2
-3.95275084E+04-8.32515675E+01-6.30156824E-03+8.01495977E-02-6.42108793E-05    3
+2.73711292E-08-4.76268611E-12-3.27129034E+04+2.84639321E+01+0.00000000E+00    4
DC5H11O2H  17/8/15      C   5H  12O   2    0G   300.000  5000.000 1397.000    61
+2.08513274E+01+2.60811030E-02-8.91735578E-06+1.38397232E-09-8.02716539E-14    2
-3.77194279E+04-8.11417120E+01-4.76374815E-01+7.83789321E-02-5.91712555E-05    3
+2.38263919E-08-3.97732270E-12-3.05087904E+04+3.26082741E+01+0.00000000E+00    4
AC5H11O2   17/8/15      C   5H  11O   2    0G   300.000  5000.000 1396.000    51
+1.98700905E+01+2.47772405E-02-8.46413614E-06+1.31283774E-09-7.61129402E-14    2
-2.04831687E+04-7.43156588E+01+3.54375282E-01+7.21758552E-02-5.35556462E-05    3
+2.12668171E-08-3.51577739E-12-1.38320365E+04+2.99444593E+01+0.00000000E+00    4
BC5H11O2   17/8/15      C   5H  11O   2    0G   300.000  5000.000 1386.000    51
+1.97546009E+01+2.47324523E-02-8.41611775E-06+1.30187335E-09-7.53316999E-14    2
-2.44671820E+04-7.68414190E+01+1.53424363E+00+6.94504944E-02-5.16917529E-05    3
+2.08690207E-08-3.52552510E-12-1.82806722E+04+2.03720098E+01+0.00000000E+00    4
CC5H11O2   17/8/15      C   5H  11O   2    0G   300.000  5000.000 1405.000    51
+2.02075561E+01+2.39554458E-02-8.06286681E-06+1.23797865E-09-7.12608001E-14    2
-2.23074093E+04-7.73358025E+01+7.15981794E-01+7.44249188E-02-5.92758872E-05    3
+2.52115515E-08-4.38572885E-12-1.60198108E+04+2.56128856E+01+0.00000000E+00    4
DC5H11O2   17/8/15      C   5H  11O   2    0G   300.000  5000.000 1396.000    51
+1.98700905E+01+2.47772405E-02-8.46413614E-06+1.31283774E-09-7.61129402E-14    2
-2.04831687E+04-7.50051405E+01+3.54375282E-01+7.21758552E-02-5.35556462E-05    3
+2.12668171E-08-3.51577739E-12-1.38320365E+04+2.92549776E+01+0.00000000E+00    4
AC5H11O    17/8/15      C   5H  11O   1    0G   300.000  5000.000 1400.000    41
+1.82339413E+01+2.37923987E-02-8.07056384E-06+1.24592855E-09-7.19996103E-14    2
-1.87450473E+04-6.87958505E+01+8.43924842E-01+6.29723769E-02-4.12079336E-05    3
+1.37396229E-08-1.84097585E-12-1.25819035E+04+2.50753974E+01+0.00000000E+00    4
BC5H11O    17/8/15      C   5H  11O   1    0G   300.000  5000.000 1378.000    41
+1.85549393E+01+2.44786662E-02-8.51926880E-06+1.33803108E-09-7.82547188E-14    2
-2.23664355E+04-7.33946136E+01+3.67366095E+00+5.17139422E-02-2.49457898E-05    3
+4.54084943E-09-3.31184982E-14-1.63228000E+04+9.40461313E+00+0.00000000E+00    4
CC5H11O    17/8/15      C   5H  11O   1    0G   300.000  5000.000 1409.000    41
+1.83213656E+01+2.35429297E-02-7.94470460E-06+1.22205357E-09-7.04356618E-14    2
-2.06340316E+04-7.05656058E+01+6.91613929E-01+6.60697133E-02-4.75285795E-05    3
+1.81072449E-08-2.84499699E-12-1.46546569E+04+2.36233979E+01+0.00000000E+00    4
DC5H11O    17/8/15      C   5H  11O   1    0G   300.000  5000.000 1400.000    41
+1.82339413E+01+2.37923987E-02-8.07056384E-06+1.24592855E-09-7.19996103E-14    2
-1.87450473E+04-6.94853322E+01+8.43924842E-01+6.29723769E-02-4.12079336E-05    3
+1.37396229E-08-1.84097585E-12-1.25819035E+04+2.43859158E+01+0.00000000E+00    4
AC5H10OOH-A 17/8/15     C   5H  11O   2    0G   300.000  5000.000 1398.000    61
+2.02759160E+01+2.40402125E-02-8.21726177E-06+1.27508622E-09-7.39470430E-14    2
-1.25890306E+04-7.45432540E+01-8.93967860E-02+7.48083410E-02-5.79088207E-05    3
+2.38676428E-08-4.05836117E-12-5.79120759E+03+3.37720278E+01+0.00000000E+00    4
AC5H10OOH-B 17/8/15     C   5H  11O   2    0G   300.000  5000.000 1390.000    61
+1.90362050E+01+2.51437855E-02-8.60836129E-06+1.33715660E-09-7.76005723E-14    2
-1.49721354E+04-6.67702235E+01+3.65133886E+00+5.70948447E-02-3.30634881E-05    3
+9.52430167E-09-1.08604128E-12-9.15524576E+03+1.73958096E+01+0.00000000E+00    4
AC5H10OOH-C 17/8/15     C   5H  11O   2    0G   300.000  5000.000 1402.000    61
+1.94269993E+01+2.45167400E-02-8.32902433E-06+1.28716724E-09-7.44370182E-14    2
-1.38808710E+04-6.93043169E+01+1.24166589E+00+6.55076365E-02-4.30153204E-05    3
+1.43717235E-08-1.92812556E-12-7.43857517E+03+2.88519661E+01+0.00000000E+00    4
AC5H10OOH-D 17/8/15     C   5H  11O   2    0G   300.000  5000.000 1398.000    61
+2.02759160E+01+2.40402125E-02-8.21726177E-06+1.27508622E-09-7.39470430E-14    2
-1.25890306E+04-7.45432540E+01-8.93967860E-02+7.48083410E-02-5.79088207E-05    3
+2.38676428E-08-4.05836117E-12-5.79120759E+03+3.37720278E+01+0.00000000E+00    4
BC5H10OOH-A 17/8/15     C   5H  11O   2    0G   300.000  5000.000 1389.000    61
+2.03178088E+01+2.39005589E-02-8.14494395E-06+1.26119353E-09-7.30298864E-14    2
-1.66270976E+04-7.71008850E+01+1.67959171E+00+7.03876561E-02-5.38977495E-05    3
+2.22634984E-08-3.82052820E-12-1.03820042E+04+2.20634050E+01+0.00000000E+00    4
BC5H10OOH-C 17/8/15     C   5H  11O   2    0G   300.000  5000.000 1390.000    61
+1.99231299E+01+2.42352995E-02-8.26025374E-06+1.27917150E-09-7.40756855E-14    2
-1.78272692E+04-7.57847609E+01+2.66396895E+00+6.53351355E-02-4.66109297E-05    3
+1.79783399E-08-2.91993271E-12-1.18409318E+04+1.67474134E+01+0.00000000E+00    4
BC5H10OOH-D 17/8/15     C   5H  11O   2    0G   300.000  5000.000 1389.000    61
+2.01548441E+01+2.39990126E-02-8.17021719E-06+1.26424565E-09-7.31718505E-14    2
-1.65704721E+04-7.70357450E+01+1.11609641E+00+7.19622376E-02-5.58678130E-05    3
+2.33617578E-08-4.04450304E-12-1.02434790E+04+2.40826139E+01+0.00000000E+00    4
CC5H10OOH-A 17/8/15     C   5H  11O   2    0G   300.000  5000.000 1407.000    61
+2.05911398E+01+2.32493648E-02-7.82909968E-06+1.20250807E-09-6.92366559E-14    2
-1.44047280E+04-7.67476901E+01+3.28493553E-01+7.68086128E-02-6.32799786E-05    3
+2.76118292E-08-4.88689574E-12-7.98741223E+03+2.98696048E+01+0.00000000E+00    4
CC5H10OOH-B 17/8/15     C   5H  11O   2    0G   300.000  5000.000 1403.000    61
+1.93820434E+01+2.43097282E-02-8.20157483E-06+1.26129144E-09-7.26836700E-14    2
-1.67969380E+04-6.98331441E+01+3.95783406E+00+5.96255587E-02-3.92210129E-05    3
+1.37408612E-08-2.01545549E-12-1.13357528E+04+1.33114157E+01+0.00000000E+00    4
CC5H10OOH-D 17/8/15     C   5H  11O   2    0G   300.000  5000.000 1407.000    61
+2.07406543E+01+2.31706906E-02-7.81225857E-06+1.20092134E-09-6.91854899E-14    2
-1.44555167E+04-7.81145448E+01+9.13421824E-01+7.51513908E-02-6.12062984E-05    3
+2.64606190E-08-4.65308639E-12-8.12947001E+03+2.63697984E+01+0.00000000E+00    4
DC5H10OOH-A 17/8/15     C   5H  11O   2    0G   300.000  5000.000 1398.000    61
+2.02759160E+01+2.40402125E-02-8.21726177E-06+1.27508622E-09-7.39470430E-14    2
-1.25890306E+04-7.45432540E+01-8.93967860E-02+7.48083410E-02-5.79088207E-05    3
+2.38676428E-08-4.05836117E-12-5.79120759E+03+3.37720278E+01+0.00000000E+00    4
DC5H10OOH-B 17/8/15     C   5H  11O   2    0G   300.000  5000.000 1390.000    61
+1.92228072E+01+2.50236156E-02-8.57782354E-06+1.33372065E-09-7.74604723E-14    2
-1.51282565E+04-6.84715050E+01+2.74458070E+00+5.78236417E-02-3.12391216E-05    3
+7.31571468E-09-4.50890257E-13-8.81862238E+03+2.20756898E+01+0.00000000E+00    4
DC5H10OOH-C 17/8/15     C   5H  11O   2    0G   300.000  5000.000 1402.000    61
+2.00395081E+01+2.42832982E-02-8.31027809E-06+1.29054421E-09-7.48846024E-14    2
-1.38460294E+04-7.39591237E+01+1.46801586E+00+6.81101661E-02-4.85321406E-05    3
+1.84083386E-08-2.91720161E-12-7.38926206E+03+2.57094934E+01+0.00000000E+00    4
A-AC5H10O  17/8/15      C   5H  10O   1    0G   300.000  5000.000 1452.000    21
+1.58864128E+01+2.27072724E-02-7.40383518E-06+1.11238546E-09-6.30611661E-14    2
-2.37201682E+04-6.09113819E+01-7.03245567E+00+8.38427156E-02-6.94901080E-05    3
+2.94315450E-08-4.93197232E-12-1.67184162E+04+5.91467747E+01+0.00000000E+00    4
A-BC5H10O  17/8/15      C   5H  10O   1    0G   300.000  5000.000 1424.000    31
+1.66888391E+01+2.23672932E-02-7.44828561E-06+1.13557959E-09-6.50516730E-14    2
-2.63127117E+04-6.48349416E+01-2.81578161E+00+7.04149950E-02-5.23593700E-05    3
+1.99929340E-08-3.05569594E-12-1.99079507E+04+3.88311343E+01+0.00000000E+00    4
A-CC5H10O  17/8/15      C   5H  10O   1    0G   300.000  5000.000 1429.000    21
+1.62176252E+01+2.18775843E-02-7.00340935E-06+1.03851279E-09-5.83155214E-14    2
-2.60452902E+04-6.25262539E+01-7.16060704E+00+8.70140494E-02-7.59660975E-05    3
+3.37198215E-08-5.87392870E-12-1.92027788E+04+5.89164749E+01+0.00000000E+00    4
A-DC5H10O  17/8/15      C   5H  10O   1    0G   300.000  5000.000 1453.000    11
+1.53604709E+01+2.35100197E-02-7.66793178E-06+1.15245719E-09-6.53534048E-14    2
-3.42487879E+04-5.88396065E+01-8.99708918E+00+8.81388493E-02-7.28825964E-05    3
+3.06897382E-08-5.10685687E-12-2.67791824E+04+6.88674277E+01+0.00000000E+00    4
B-CC5H10O  9/ 8/14      C   5H  10O   1    0G   300.000  5000.000 1413.000    31
+1.72822083E+01+2.21811831E-02-7.45086135E-06+1.14266526E-09-6.57264262E-14    2
-2.89756909E+04-6.99425869E+01-4.02733813E+00+7.75766076E-02-6.31068363E-05    3
+2.66344724E-08-4.52085229E-12-2.22133168E+04+4.23801047E+01+0.00000000E+00    4
B-DC5H10O  9/ 8/14      C   5H  10O   1    0G   300.000  5000.000 1426.000    21
+1.59398262E+01+2.34035968E-02-7.80111462E-06+1.19023227E-09-6.82188270E-14    2
-2.75659851E+04-6.31518634E+01-4.57207704E+00+7.33362569E-02-5.36913946E-05    3
+2.00360735E-08-2.97590047E-12-2.07808158E+04+4.60627306E+01+0.00000000E+00    4
C-DC5H10O  17/8/15      C   5H  10O   1    0G   300.000  5000.000 1415.000    31
+1.75721707E+01+2.16805796E-02-7.22379193E-06+1.10170103E-09-6.31222440E-14    2
-2.54336652E+04-7.01131722E+01-7.94334743E+00+9.36350437E-02-8.55713608E-05    3
+3.97013264E-08-7.24456558E-12-1.79116899E+04+6.23627456E+01+0.00000000E+00    4
AC5H10OOH-AO2 8/15      C   5H  11O   4    0G   300.000  5000.000 1397.000    71
+2.49284926E+01+2.49502228E-02-8.57455029E-06+1.33547829E-09-7.76537998E-14    2
-3.17167911E+04-9.46333090E+01+1.47959220E+00+8.37668710E-02-6.63705552E-05    3
+2.76480297E-08-4.71460623E-12-2.39474084E+04+2.99187562E+01+0.00000000E+00    4
AC5H10OOH-BO2 8/15      C   5H  11O   4    0G   300.000  5000.000 1389.000    71
+2.48032671E+01+2.49329192E-02-8.54000436E-06+1.32701219E-09-7.70333881E-14    2
-3.56964132E+04-9.64200661E+01+2.66224628E+00+8.10932443E-02-6.46324438E-05    3
+2.73538724E-08-4.75157092E-12-2.83982547E+04+2.10041880E+01+0.00000000E+00    4
AC5H10OOH-CO2 8/15      C   5H  11O   4    0G   300.000  5000.000 1405.000    71
+2.52420639E+01+2.41694359E-02-8.19141254E-06+1.26381882E-09-7.30015120E-14    2
-3.35305240E+04-9.68327377E+01+1.83495697E+00+8.60948213E-02-7.22651143E-05    3
+3.17312304E-08-5.62009843E-12-2.61355447E+04+2.62902691E+01+0.00000000E+00    4
AC5H10OOH-DO2 8/15      C   5H  11O   4    0G   300.000  5000.000 1397.000    71
+2.49284926E+01+2.49502228E-02-8.57455029E-06+1.33547829E-09-7.76537998E-14    2
-3.17167911E+04-9.46333090E+01+1.47959220E+00+8.37668710E-02-6.63705552E-05    3
+2.76480297E-08-4.71460623E-12-2.39474084E+04+2.99187562E+01+0.00000000E+00    4
BC5H10OOH-AO2 8/15      C   5H  11O   4    0G   300.000  5000.000 1389.000    71
+2.48032671E+01+2.49329192E-02-8.54000436E-06+1.32701219E-09-7.70333881E-14    2
-3.56964132E+04-9.64200661E+01+2.66224628E+00+8.10932443E-02-6.46324438E-05    3
+2.73538724E-08-4.75157092E-12-2.83982547E+04+2.10041880E+01+0.00000000E+00    4
BC5H10OOH-CO2 8/15      C   5H  11O   4    0G   300.000  5000.000 1396.000    71
+2.51614268E+01+2.40667268E-02-8.11773937E-06+1.24830451E-09-7.19346846E-14    2
-3.75274060E+04-9.95533661E+01+2.92757922E+00+8.37497935E-02-7.09476834E-05    3
+3.16521003E-08-5.69638239E-12-3.05708429E+04+1.71231211E+01+0.00000000E+00    4
BC5H10OOH-DO2 8/15      C   5H  11O   4    0G   300.000  5000.000 1389.000    71
+2.48032671E+01+2.49329192E-02-8.54000436E-06+1.32701219E-09-7.70333881E-14    2
-3.56964132E+04-9.71095477E+01+2.66224628E+00+8.10932443E-02-6.46324438E-05    3
+2.73538724E-08-4.75157092E-12-2.83982547E+04+2.03147064E+01+0.00000000E+00    4
CC5H10OOH-AO2 8/15      C   5H  11O   4    0G   300.000  5000.000 1405.000    71
+2.52420639E+01+2.41694359E-02-8.19141254E-06+1.26381882E-09-7.30015120E-14    2
-3.35305240E+04-9.68327377E+01+1.83495697E+00+8.60948213E-02-7.22651143E-05    3
+3.17312304E-08-5.62009843E-12-2.61355447E+04+2.62902691E+01+0.00000000E+00    4
CC5H10OOH-BO2 8/15      C   5H  11O   4    0G   300.000  5000.000 1396.000    71
+2.51614268E+01+2.40667268E-02-8.11773937E-06+1.24830451E-09-7.19346846E-14    2
-3.75274060E+04-9.95533661E+01+2.92757922E+00+8.37497935E-02-7.09476834E-05    3
+3.16521003E-08-5.69638239E-12-3.05708429E+04+1.71231211E+01+0.00000000E+00    4
CC5H10OOH-DO2 8/15      C   5H  11O   4    0G   300.000  5000.000 1405.000    71
+2.52420639E+01+2.41694359E-02-8.19141254E-06+1.26381882E-09-7.30015120E-14    2
-3.35305240E+04-9.75222193E+01+1.83495697E+00+8.60948213E-02-7.22651143E-05    3
+3.17312304E-08-5.62009843E-12-2.61355447E+04+2.56007875E+01+0.00000000E+00    4
DC5H10OOH-AO2 8/15      C   5H  11O   4    0G   300.000  5000.000 1397.000    71
+2.49284926E+01+2.49502228E-02-8.57455029E-06+1.33547829E-09-7.76537998E-14    2
-3.17167911E+04-9.46333090E+01+1.47959220E+00+8.37668710E-02-6.63705552E-05    3
+2.76480297E-08-4.71460623E-12-2.39474084E+04+2.99187562E+01+0.00000000E+00    4
DC5H10OOH-BO2 8/15      C   5H  11O   4    0G   300.000  5000.000 1389.000    71
+2.48032671E+01+2.49329192E-02-8.54000436E-06+1.32701219E-09-7.70333881E-14    2
-3.56964132E+04-9.71095477E+01+2.66224628E+00+8.10932443E-02-6.46324438E-05    3
+2.73538724E-08-4.75157092E-12-2.83982547E+04+2.03147064E+01+0.00000000E+00    4
DC5H10OOH-CO2 8/15      C   5H  11O   4    0G   300.000  5000.000 1405.000    71
+2.52420639E+01+2.41694359E-02-8.19141254E-06+1.26381882E-09-7.30015120E-14    2
-3.35305240E+04-9.75222193E+01+1.83495697E+00+8.60948213E-02-7.22651143E-05    3
+3.17312304E-08-5.62009843E-12-2.61355447E+04+2.56007875E+01+0.00000000E+00    4
C5H9A-A,BOOH  8/15      C   5H  11O   4    0G   300.000  5000.000 1391.000    81
+2.53148126E+01+2.41050499E-02-8.26152052E-06+1.28429464E-09-7.45769254E-14    2
-2.78251062E+04-9.70436295E+01+2.87832948E+00+8.17084683E-02-6.64693824E-05    3
+2.85545390E-08-5.00710723E-12-2.05092635E+04+2.16842979E+01+0.00000000E+00    4
C5H9A-A,COOH  8/15      C   5H  11O   4    0G   300.000  5000.000 1406.000    81
+2.55933245E+01+2.34677500E-02-7.95418684E-06+1.22729993E-09-7.08960495E-14    2
-2.56096120E+04-9.67335324E+01+1.46543304E+00+8.83867154E-02-7.62009797E-05    3
+3.41128921E-08-6.11972135E-12-1.81049887E+04+2.97796524E+01+0.00000000E+00    4
C5H9A-A,DOOH  8/15      C   5H  11O   4    0G   300.000  5000.000 1399.000    81
+2.53362233E+01+2.42043007E-02-8.32306052E-06+1.29685010E-09-7.54306895E-14    2
-2.38227509E+04-9.48747338E+01+1.03378269E+00+8.63930746E-02-7.07031565E-05    3
+3.02282342E-08-5.25110249E-12-1.59058366E+04+3.37540294E+01+0.00000000E+00    4
C5H9A-B,COOH  8/15      C   5H  11O   4    0G   300.000  5000.000 1398.000    81
+2.56997668E+01+2.32725079E-02-7.86284471E-06+1.21047841E-09-6.98107824E-14    2
-2.96771591E+04-9.96712347E+01+3.12194965E+00+8.44868328E-02-7.28869575E-05    3
+3.29012852E-08-5.96274974E-12-2.26799790E+04+1.85842452E+01+0.00000000E+00    4
C5H9A-B,DOOH  8/15      C   5H  11O   4    0G   300.000  5000.000 1391.000    81
+2.53148126E+01+2.41050499E-02-8.26152052E-06+1.28429464E-09-7.45769254E-14    2
-2.78251062E+04-9.70436295E+01+2.87832948E+00+8.17084683E-02-6.64693824E-05    3
+2.85545390E-08-5.00710723E-12-2.05092635E+04+2.16842979E+01+0.00000000E+00    4
C5H9A-C,DOOH  8/15      C   5H  11O   4    0G   300.000  5000.000 1406.000    81
+2.55933245E+01+2.34677500E-02-7.95418684E-06+1.22729993E-09-7.08960495E-14    2
-2.56096120E+04-9.67335324E+01+1.46543304E+00+8.83867154E-02-7.62009797E-05    3
+3.41128921E-08-6.11972135E-12-1.81049887E+04+2.97796524E+01+0.00000000E+00    4
C5H9B-A,AOOH  8/15      C   5H  11O   4    0G   300.000  5000.000 1392.000    81
+2.37032599E+01+2.57553915E-02-8.89408554E-06+1.38970172E-09-8.09866916E-14    2
-2.62015201E+04-8.58515282E+01+4.28350134E+00+6.83511301E-02-4.42293137E-05    3
+1.46614813E-08-1.99882623E-12-1.91209818E+04+1.95267791E+01+0.00000000E+00    4
C5H9B-A,COOH  8/15      C   5H  11O   4    0G   300.000  5000.000 1675.000    81
+2.44195505E+01+2.45182960E-02-8.32768546E-06+1.28669810E-09-7.43971425E-14    2
-2.80210816E+04-8.93466817E+01+5.06775026E+00+7.13339940E-02-5.22649130E-05    3
+2.02919064E-08-3.25625167E-12-2.14500744E+04+1.40310906E+01+0.00000000E+00    4
C5H9B-A,DOOH  8/15      C   5H  11O   4    0G   300.000  5000.000 1392.000    81
+2.37032599E+01+2.57553915E-02-8.89408554E-06+1.38970172E-09-8.09866916E-14    2
-2.62015201E+04-8.51620466E+01+4.28350134E+00+6.83511301E-02-4.42293137E-05    3
+1.46614813E-08-1.99882623E-12-1.91209818E+04+2.02162608E+01+0.00000000E+00    4
C5H9B-C,DOOH  8/15      C   5H  11O   4    0G   300.000  5000.000 1675.000    81
+2.44195505E+01+2.45182960E-02-8.32768546E-06+1.28669810E-09-7.43971425E-14    2
-2.80210816E+04-9.07256450E+01+5.06775026E+00+7.13339940E-02-5.22649130E-05    3
+2.02919064E-08-3.25625167E-12-2.14500744E+04+1.26521274E+01+0.00000000E+00    4
C5H9C-A,AOOH  8/15      C   5H  11O   4    0G   300.000  5000.000 1681.000    81
+2.63011187E+01+2.38231644E-02-8.29527214E-06+1.30384489E-09-7.63133641E-14    2
-2.62801782E+04-1.01764259E+02+2.40737385E+00+7.31844750E-02-4.34551328E-05    3
+1.06843813E-08-6.06073375E-13-1.74826725E+04+2.86070302E+01+0.00000000E+00    4
C5H9C-A,BOOH  8/15      C   5H  11O   4    0G   300.000  5000.000 1393.000    81
+2.49289305E+01+2.44398284E-02-8.37848298E-06+1.30269965E-09-7.56543783E-14    2
-2.90312299E+04-9.50950095E+01+3.83902707E+00+7.67534526E-02-5.93019661E-05    3
+2.43350243E-08-4.12011052E-12-2.19645331E+04+1.71683879E+01+0.00000000E+00    4
C5H9C-A,DOOH  8/15      C   5H  11O   4    0G   300.000  5000.000 1681.000    81
+2.63011187E+01+2.38231644E-02-8.29527214E-06+1.30384489E-09-7.63133641E-14    2
-2.62801782E+04-1.01074777E+02+2.40737385E+00+7.31844750E-02-4.34551328E-05    3
+1.06843813E-08-6.06073375E-13-1.74826725E+04+2.92965119E+01+0.00000000E+00    4
C5H9C-B,DOOH  8/15      C   5H  11O   4    0G   300.000  5000.000 1393.000    81
+2.49289305E+01+2.44398284E-02-8.37848298E-06+1.30269965E-09-7.56543783E-14    2
-2.90312299E+04-9.57844912E+01+3.83902707E+00+7.67534526E-02-5.93019661E-05    3
+2.43350243E-08-4.12011052E-12-2.19645331E+04+1.64789063E+01+0.00000000E+00    4
C5H9D-A,AOOH  8/15      C   5H  11O   4    0G   300.000  5000.000 1399.000    81
+2.53362233E+01+2.42043007E-02-8.32306052E-06+1.29685010E-09-7.54306895E-14    2
-2.38227509E+04-9.55642154E+01+1.03378269E+00+8.63930746E-02-7.07031565E-05    3
+3.02282342E-08-5.25110249E-12-1.59058366E+04+3.30645478E+01+0.00000000E+00    4
C5H9D-A,BOOH  8/15      C   5H  11O   4    0G   300.000  5000.000 1391.000    81
+2.51743725E+01+2.42094413E-02-8.29427020E-06+1.28906994E-09-7.48414448E-14    2
-2.77836927E+04-9.64353283E+01+2.27985031E+00+8.34372048E-02-6.86098141E-05    3
+2.97415611E-08-5.24930633E-12-2.03658212E+04+2.45531752E+01+0.00000000E+00    4
C5H9D-A,COOH  8/15      C   5H  11O   4    0G   300.000  5000.000 1406.000    81
+2.56538280E+01+2.34057032E-02-7.93032646E-06+1.22331141E-09-7.06528620E-14    2
-2.56105413E+04-9.68592428E+01+2.13973267E+00+8.63107772E-02-7.36971527E-05    3
+3.27651712E-08-5.85073945E-12-1.82585105E+04+2.65675140E+01+0.00000000E+00    4
C5H9D-B,COOH  8/15      C   5H  11O   4    0G   300.000  5000.000 1398.000    81
+2.56997668E+01+2.32725079E-02-7.86284471E-06+1.21047841E-09-6.98107824E-14    2
-2.96771591E+04-1.00360716E+02+3.12194965E+00+8.44868328E-02-7.28869575E-05    3
+3.29012852E-08-5.96274974E-12-2.26799790E+04+1.78947636E+01+0.00000000E+00    4
C5H9A-AOOH 9/ 8/14      C   5H  10O   2    0G   300.000  5000.000 1388.000    51
+2.12338541E+01+2.14695668E-02-7.41711017E-06+1.15964346E-09-6.76214281E-14    2
-2.22824726E+04-8.15535062E+01-5.66437031E-01+7.51592771E-02-5.92588303E-05    3
+2.44464873E-08-4.14011509E-12-1.49441419E+04+3.46236211E+01+0.00000000E+00    4
C5H9A-COOH 9/ 8/14      C   5H  10O   2    0G   300.000  5000.000 1396.000    51
+2.21762503E+01+2.02997794E-02-6.93527858E-06+1.07653985E-09-6.24712973E-14    2
-2.45061123E+04-8.96059444E+01-2.23218718E+00+8.31068782E-02-6.96695008E-05    3
+2.98090622E-08-5.11291423E-12-1.66665651E+04+3.93336979E+01+0.00000000E+00    4
C5H9A-DOOH 9/ 8/14      C   5H  10O   2    0G   300.000  5000.000 1393.000    51
+1.91192483E+01+2.31083713E-02-7.94263265E-06+1.23713692E-09-7.19377465E-14    2
-2.31563003E+04-7.06976781E+01+5.84051402E-01+6.61435369E-02-4.64794214E-05    3
+1.71320929E-08-2.62129070E-12-1.66564666E+04+2.90021482E+01+0.00000000E+00    4
C5H9B-AOOH 9/ 8/14      C   5H  10O   2    0G   300.000  5000.000 1385.000    51
+2.11330268E+01+2.15086873E-02-7.42113144E-06+1.15934717E-09-6.75687044E-14    2
-2.35608139E+04-8.15040563E+01+5.49656384E-01+7.04990310E-02-5.27825801E-05    3
+2.06470792E-08-3.33664189E-12-1.64635942E+04+2.87891957E+01+0.00000000E+00    4
C5H9B-DOOH 9/ 8/14      C   5H  10O   2    0G   300.000  5000.000 1385.000    51
+2.11330268E+01+2.15086873E-02-7.42113144E-06+1.15934717E-09-6.75687044E-14    2
-2.35608139E+04-8.15040563E+01+5.49656384E-01+7.04990310E-02-5.27825801E-05    3
+2.06470792E-08-3.33664189E-12-1.64635942E+04+2.87891957E+01+0.00000000E+00    4
C5H9C-AOOH 9/ 8/14      C   5H  10O   2    0G   300.000  5000.000 1396.000    51
+1.95116301E+01+2.27723060E-02-7.82629606E-06+1.21895173E-09-7.08783753E-14    2
-2.27377278E+04-7.28224624E+01-1.33187657E-02+6.92568397E-02-5.06647207E-05    3
+1.94153559E-08-3.06921462E-12-1.60254301E+04+3.17599798E+01+0.00000000E+00    4
C5H9C-BOOH 9/ 8/14      C   5H  10O   2    0G   300.000  5000.000 1393.000    51
+2.30088665E+01+1.91355851E-02-6.44358123E-06+9.91225120E-10-5.71817398E-14    2
-2.66103173E+04-9.24108219E+01-1.04862343E+00+8.26699722E-02-7.17941940E-05    3
+3.18245309E-08-5.62912876E-12-1.90383401E+04+3.41116802E+01+0.00000000E+00    4
C5H9OA-AOOH-B 8/15      C   5H  10O   3    0G   300.000  5000.000 1421.000    41
+2.17927261E+01+2.30720633E-02-7.77386468E-06+1.19507605E-09-6.88699665E-14    2
-3.96712246E+04-8.94813847E+01-5.49708925E+00+9.47288852E-02-8.00296268E-05    3
+3.42124943E-08-5.80022917E-12-3.11441575E+04+5.40078635E+01+0.00000000E+00    4
C5H9OA-AOOH-C 8/15      C   5H  10O   3    0G   300.000  5000.000 1426.000    41
+2.27244179E+01+2.20779072E-02-7.39099655E-06+1.13153303E-09-6.50287263E-14    2
-3.78217375E+04-9.29947975E+01-6.41150803E+00+9.94317564E-02-8.58615548E-05    3
+3.70273302E-08-6.27783473E-12-2.88551995E+04+5.98124271E+01+0.00000000E+00    4
C5H9OA-AOOH-D 8/15      C   5H  10O   3    0G   300.000  5000.000 1411.000    41
+2.16522955E+01+2.34455715E-02-7.95666190E-06+1.22905457E-09-7.10634551E-14    2
-3.55963177E+04-8.69264178E+01-8.39507263E+00+1.05102811E-01-9.37685656E-05    3
+4.22174145E-08-7.50607159E-12-2.64325286E+04+7.01690143E+01+0.00000000E+00    4
C5H9OA-BOOH-A 8/15      C   5H  10O   3    0G   300.000  5000.000 1417.000    51
+2.17022735E+01+2.26119914E-02-7.58981668E-06+1.16366327E-09-6.69308130E-14    2
-3.75365241E+04-8.49179287E+01-1.90416408E+00+8.28866784E-02-6.64998506E-05    3
+2.72221761E-08-4.44711330E-12-2.99886544E+04+3.98116691E+01+0.00000000E+00    4
C5H9OA-BOOH-C 8/15      C   5H  10O   3    0G   300.000  5000.000 1417.000    51
+2.32822727E+01+2.16339746E-02-7.33435063E-06+1.13242966E-09-6.54655290E-14    2
-4.01984498E+04-9.51976254E+01-4.48273125E-01+7.90873425E-02-5.97079860E-05    3
+2.24183926E-08-3.31048774E-12-3.23280594E+04+3.12502863E+01+0.00000000E+00    4
C5H9OA-BOOH-D 8/15      C   5H  10O   3    0G   300.000  5000.000 1417.000    51
+2.17022735E+01+2.26119914E-02-7.58981668E-06+1.16366327E-09-6.69308130E-14    2
-3.75365241E+04-8.49179287E+01-1.90416408E+00+8.28866784E-02-6.64998506E-05    3
+2.72221761E-08-4.44711330E-12-2.99886544E+04+3.98116691E+01+0.00000000E+00    4
C5H9OA-COOH-A 8/15      C   5H  10O   3    0G   300.000  5000.000 1416.000    41
+2.19787258E+01+2.27762232E-02-7.64127053E-06+1.17119291E-09-6.73502124E-14    2
-3.79400480E+04-8.78800726E+01-8.23567336E+00+1.06958451E-01-9.80175480E-05    3
+4.50653157E-08-8.12667607E-12-2.89611267E+04+6.93052953E+01+0.00000000E+00    4
C5H9OA-COOH-B 8/15      C   5H  10O   3    0G   300.000  5000.000 1427.000    41
+2.18581268E+01+2.26582661E-02-7.55183274E-06+1.15215111E-09-6.60356238E-14    2
-4.18939906E+04-8.96205075E+01-6.82291569E+00+1.03424198E-01-9.51789693E-05    3
+4.41170689E-08-8.01854503E-12-3.34508247E+04+5.92928651E+01+0.00000000E+00    4
C5H9OA-COOH-D 8/15      C   5H  10O   3    0G   300.000  5000.000 1416.000    41
+2.19787258E+01+2.27762232E-02-7.64127053E-06+1.17119291E-09-6.73502124E-14    2
-3.79400480E+04-8.78800726E+01-8.23567336E+00+1.06958451E-01-9.80175480E-05    3
+4.50653157E-08-8.12667607E-12-2.89611267E+04+6.93052953E+01+0.00000000E+00    4
C5H9OA-DOOH-A 8/15      C   5H  10O   3    0G   300.000  5000.000 1412.000    31
+2.10306351E+01+2.43651936E-02-8.26752696E-06+1.27699187E-09-7.38333381E-14    2
-4.61055228E+04-8.36588979E+01-1.05445809E+01+1.09794719E-01-9.75108462E-05    3
+4.36190126E-08-7.70228936E-12-3.64529482E+04+8.15338458E+01+0.00000000E+00    4
C5H9OA-DOOH-B 8/15      C   5H  10O   3    0G   300.000  5000.000 1424.000    31
+2.09160528E+01+2.42617893E-02-8.18691855E-06+1.25968394E-09-7.26328496E-14    2
-5.00500176E+04-8.54043566E+01-8.94627226E+00+1.05725319E-01-9.40624065E-05    3
+4.23682039E-08-7.53895269E-12-4.09789989E+04+7.06042654E+01+0.00000000E+00    4
C5H9OA-DOOH-C 8/15      C   5H  10O   3    0G   300.000  5000.000 1418.000    31
+2.17931949E+01+2.35822973E-02-7.96856856E-06+1.22739410E-09-7.08291072E-14    2
-4.82483390E+04-8.87831309E+01-1.00859009E+01+1.11154142E-01-1.00718064E-04    3
+4.57405620E-08-8.16324506E-12-3.86489157E+04+7.75075179E+01+0.00000000E+00    4
C5H9OB-COOH-A 8/15      C   5H  10O   3    0G   300.000  5000.000 1427.000    51
+2.33660026E+01+2.12967547E-02-7.16311642E-06+1.10028483E-09-6.33839052E-14    2
-4.02710909E+04-9.55650042E+01-2.03626914E+00+8.44316222E-02-6.63448448E-05    3
+2.58620472E-08-3.95367034E-12-3.20450331E+04+3.91516619E+01+0.00000000E+00    4
C5H9OB-COOH-D 8/15      C   5H  10O   3    0G   300.000  5000.000 1427.000    51
+2.33660026E+01+2.12967547E-02-7.16311642E-06+1.10028483E-09-6.33839052E-14    2
-4.02710909E+04-9.62544859E+01-2.03626914E+00+8.44316222E-02-6.63448448E-05    3
+2.58620472E-08-3.95367034E-12-3.20450331E+04+3.84621803E+01+0.00000000E+00    4
C5H9OB-DOOH-A 9/14      C   5H  10O   3    0G   300.000  5000.000 1420.000    41
+2.09989877E+01+2.35749161E-02-7.91024357E-06+1.21256198E-09-6.97360491E-14    2
-3.87964686E+04-8.27787933E+01-3.52560638E+00+8.53243101E-02-6.71300274E-05    3
+2.68114187E-08-4.26214321E-12-3.08855835E+04+4.70812100E+01+0.00000000E+00    4
C5H9OB-DOOH-C 9/14      C   5H  10O   3    0G   300.000  5000.000 1416.000    41
+2.23010712E+01+2.28353062E-02-7.73563047E-06+1.19365671E-09-6.89722094E-14    2
-4.13407064E+04-9.21482846E+01-3.01430534E+00+8.55622233E-02-6.67458085E-05    3
+2.61563238E-08-4.06382943E-12-3.30739466E+04+4.22585328E+01+0.00000000E+00    4
C5H9OC-DOOH-A 8/15      C   5H  10O   3    0G   300.000  5000.000 1424.000    51
+2.32181188E+01+2.12380409E-02-7.10087806E-06+1.08610144E-09-6.23742333E-14    2
-3.68812122E+04-9.30381675E+01-4.71787956E+00+9.63722654E-02-8.44994419E-05    3
+3.70849590E-08-6.39906257E-12-2.83656016E+04+5.31581269E+01+0.00000000E+00    4
C5H9OC-DOOH-B 8/15      C   5H  10O   3    0G   300.000  5000.000 1424.000    51
+2.31592020E+01+2.11055768E-02-7.01494893E-06+1.06850406E-09-6.11803452E-14    2
-4.08758474E+04-9.58608672E+01-3.31967698E+00+9.28312807E-02-8.14721652E-05    3
+3.59633071E-08-6.24713097E-12-3.28520059E+04+4.25342095E+01+0.00000000E+00    4
CH3COCH2OCH2CH2 14      C   5H   9O   2    0G   300.000  5000.000 1398.000    51
+1.61915801E+01+2.17259962E-02-7.18255818E-06+1.08967551E-09-6.22058703E-14    2
-2.83312411E+04-5.06778787E+01+2.46265398E+00+5.31605978E-02-3.44158813E-05    3
+1.17106545E-08-1.63587278E-12-2.35149168E+04+2.32544951E+01+0.00000000E+00    4
IC5KETAA   17/8/15      C   5H  10O   3    0G   300.000  5000.000 1396.000    61
+2.14062122E+01+2.31814714E-02-7.94585296E-06+1.23549697E-09-7.17602293E-14    2
-4.77416322E+04-7.94699242E+01+2.55453432E+00+6.48725206E-02-4.21449634E-05    3
+1.35396181E-08-1.69771989E-12-4.09936393E+04+2.25509833E+01+0.00000000E+00    4
IC5KETAB   17/8/15      C   5H  10O   3    0G   300.000  5000.000 1387.000    61
+2.54563544E+01+2.01871439E-02-7.02056943E-06+1.10298380E-09-6.45487927E-14    2
-5.08666110E+04-1.03884759E+02-2.76644890E-01+8.19422293E-02-6.36165752E-05    3
+2.46645924E-08-3.82375149E-12-4.21788557E+04+3.35972645E+01+0.00000000E+00    4
IC5KETAC   17/8/15      C   5H  10O   3    0G   300.000  5000.000 1530.000    61
+2.36202007E+01+2.16574723E-02-7.50493626E-06+1.17597427E-09-6.86855912E-14    2
-5.08399014E+04-9.37964825E+01+3.38364660E+00+6.08702747E-02-3.15372777E-05    3
+4.94036887E-09+4.82022927E-13-4.31638560E+04+1.74830999E+01+0.00000000E+00    4
IC5KETAD   17/8/15      C   5H  10O   3    0G   300.000  5000.000 1396.000    61
+2.14062122E+01+2.31814714E-02-7.94585296E-06+1.23549697E-09-7.17602293E-14    2
-4.77416322E+04-7.94699242E+01+2.55453432E+00+6.48725206E-02-4.21449634E-05    3
+1.35396181E-08-1.69771989E-12-4.09936393E+04+2.25509833E+01+0.00000000E+00    4
IC5KETCA   17/8/15      C   5H  10O   3    0G   300.000  5000.000 1403.000    61
+1.99169154E+01+2.37975805E-02-8.01511093E-06+1.23140060E-09-7.09187874E-14    2
-5.11169360E+04-7.05780003E+01+3.30504848E+00+6.12212470E-02-3.95733068E-05    3
+1.30417749E-08-1.72022312E-12-4.52388966E+04+1.90774795E+01+0.00000000E+00    4
IC5KETCB   17/8/15      C   5H  10O   3    0G   300.000  5000.000 1388.000    61
+2.43081284E+01+2.03116947E-02-6.88557448E-06+1.06413626E-09-6.15901378E-14    2
-5.43890101E+04-9.76241400E+01+4.99341353E-01+7.79929244E-02-6.02225926E-05    3
+2.34360987E-08-3.65044242E-12-4.64243747E+04+2.93525587E+01+0.00000000E+00    4
IC5KETCD   17/8/15      C   5H  10O   3    0G   300.000  5000.000 1394.000    61
+2.37898908E+01+2.04031709E-02-6.84168010E-06+1.04954951E-09-6.04313994E-14    2
-5.08956742E+04-9.25390969E+01-2.83543507E-01+8.06299025E-02-6.46191514E-05    3
+2.62468255E-08-4.26140982E-12-4.30486170E+04+3.51463538E+01+0.00000000E+00    4
IC5KETDA   17/8/15      C   5H  10O   3    0G   300.000  5000.000 1395.000    61
+2.23252658E+01+2.23009872E-02-7.62390887E-06+1.18364958E-09-6.86862585E-14    2
-4.79954210E+04-8.50606082E+01+1.31890291E+00+7.08408070E-02-4.98675222E-05    3
+1.76320223E-08-2.48535036E-12-4.07142424E+04+2.78334474E+01+0.00000000E+00    4
IC5KETDB   17/8/15      C   5H  10O   3    0G   300.000  5000.000 1381.000    61
+2.22545164E+01+2.21858094E-02-7.54539826E-06+1.16735178E-09-6.75734913E-14    2
-5.19970461E+04-8.78431657E+01+2.45036196E+00+6.83213847E-02-4.82822981E-05    3
+1.73840001E-08-2.52418883E-12-4.51554184E+04+1.84815016E+01+0.00000000E+00    4
IC5KETDC   17/8/15      C   5H  10O   3    0G   300.000  5000.000 1391.000    61
+2.57459735E+01+1.95157132E-02-6.70259887E-06+1.04493380E-09-6.08454008E-14    2
-4.96555982E+04-1.04885682E+02-2.47013912E+00+9.30872396E-02-8.13203099E-05    3
+3.57768012E-08-6.26400503E-12-4.06868372E+04+4.38329357E+01+0.00000000E+00    4
IC5KETAAO  17/8/15      C   5H   9O   2    0G   300.000  5000.000 1670.000    41
+1.54491093E+01+2.58830088E-02-9.38194545E-06+1.51919963E-09-9.08764412E-14    2
-2.73128942E+04-4.89349130E+01+6.20340512E+00+3.78488938E-02-8.21632367E-06    3
-4.45998794E-09+1.69104440E-12-2.33706795E+04+3.88282175E+00+0.00000000E+00    4
IC5KETABO  17/8/15      C   5H   9O   2    0G   300.000  5000.000 1680.000    41
+1.74003757E+01+2.43634015E-02-8.89217693E-06+1.44672950E-09-8.68336325E-14    2
-2.96359315E+04-6.26150618E+01+2.44492593E+00+5.39988220E-02-2.76353434E-05    3
+5.14986988E-09-2.28548561E-14-2.42538749E+04+1.91347808E+01+0.00000000E+00    4
IC5KETACO  17/8/15      C   5H   9O   2    0G   300.000  5000.000 1405.000    41
+1.87759820E+01+2.09363794E-02-7.11851372E-06+1.10072541E-09-6.36812526E-14    2
-3.10560920E+04-6.84256552E+01+3.17102493E+00+5.52252992E-02-3.48045866E-05    3
+1.07470812E-08-1.26264879E-12-2.54634549E+04+1.60763592E+01+0.00000000E+00    4
IC5KETADO  17/8/15      C   5H   9O   2    0G   300.000  5000.000 1670.000    41
+1.54491093E+01+2.58830088E-02-9.38194545E-06+1.51919963E-09-9.08764412E-14    2
-2.73128942E+04-4.89349130E+01+6.20340512E+00+3.78488938E-02-8.21632367E-06    3
-4.45998794E-09+1.69104440E-12-2.33706795E+04+3.88282175E+00+0.00000000E+00    4
IC5KETCAO  17/8/15      C   5H   9O   2    0G   300.000  5000.000 1514.000    41
+1.72485932E+01+2.16326796E-02-7.22890702E-06+1.10467817E-09-6.33813429E-14    2
-3.21371394E+04-5.86643290E+01+4.75737279E+00+4.52905574E-02-2.09520730E-05    3
+2.65371883E-09+4.60703138E-13-2.73333149E+04+1.02325004E+01+0.00000000E+00    4
IC5KETCBO  17/8/15      C   5H   9O   2    0G   300.000  5000.000 1510.000    41
+1.93742496E+01+2.06425485E-02-7.06983683E-06+1.09902869E-09-6.38342204E-14    2
-3.47003768E+04-7.43848166E+01+4.60922258E+00+4.63105317E-02-1.85546802E-05    3
-2.86158793E-10+1.27532426E-12-2.87895902E+04+7.87701574E+00+0.00000000E+00    4
IC5KETCDO  17/8/15      C   5H   9O   2    0G   300.000  5000.000 1489.000    41
+1.78986194E+01+2.13374499E-02-7.19313241E-06+1.10668165E-09-6.38266549E-14    2
-3.16063716E+04-6.33320448E+01+7.66113508E+00+3.31212888E-02-2.76253288E-06    3
-8.32131128E-09+2.78275744E-12-2.68823428E+04-4.11946991E+00+0.00000000E+00    4
IC5KETDAO  17/8/15      C   5H   9O   2    0G   300.000  5000.000 1485.000    41
+1.95835650E+01+2.02788959E-02-6.90312559E-06+1.06869517E-09-6.18931202E-14    2
-2.89934666E+04-7.27514739E+01+2.77854914E+00+5.49042648E-02-3.12957279E-05    3
+7.33340136E-09-3.35699979E-13-2.28103088E+04+1.89499650E+01+0.00000000E+00    4
IC5KETDBO  17/8/15      C   5H   9O   2    0G   300.000  5000.000 1519.000    41
+2.00669200E+01+2.02402238E-02-6.97500713E-06+1.08902290E-09-6.34524956E-14    2
-3.25858999E+04-7.80517736E+01+5.21028340E+00+4.44018385E-02-1.51327339E-05    3
-2.59536762E-09+1.79445594E-12-2.64639770E+04+5.32661738E+00+0.00000000E+00    4
IC5KETDCO  17/8/15      C   5H   9O   2    0G   300.000  5000.000 1385.000    41
+2.06749614E+01+2.01791491E-02-7.04935407E-06+1.11015087E-09-6.50552099E-14    2
-3.08738095E+04-8.00272702E+01+1.74667514E+00+6.15641942E-02-4.06488995E-05    3
+1.31250854E-08-1.65755406E-12-2.40252952E+04+2.26218438E+01+0.00000000E+00    4
AC5H10OH   17/8/15      C   5H  11O   1    0G   300.000  5000.000 1396.000    51
+1.64350382E+01+2.48732260E-02-8.43959366E-06+1.30322470E-09-7.53261177E-14    2
-2.28956938E+04-5.51681478E+01+1.23496772E+00+5.48298602E-02-2.85379159E-05    3
+6.14801654E-09-2.41162327E-13-1.70643706E+04+2.84296007E+01+0.00000000E+00    4
BC5H10OH   17/8/15      C   5H  11O   1    0G   300.000  5000.000 1384.000    51
+1.69551854E+01+2.50397308E-02-8.62897621E-06+1.34632322E-09-7.83770200E-14    2
-2.52556374E+04-6.12549178E+01+2.16094248E+00+5.26897228E-02-2.56800949E-05    3
+4.72180512E-09-1.32098054E-14-1.93564411E+04+2.07680728E+01+0.00000000E+00    4
CC5H10OH   17/8/15      C   5H  11O   1    0G   300.000  5000.000 1408.000    51
+1.76376123E+01+2.33184854E-02-7.78464125E-06+1.18857749E-09-6.81463457E-14    2
-2.21964329E+04-6.38737345E+01-1.66278849E+00+7.47656913E-02-6.14804272E-05    3
+2.69357912E-08-4.78920793E-12-1.61297989E+04+3.75225406E+01+0.00000000E+00    4
AO2C5H10OH 17/8/15      C   5H  11O   3    0G   300.000  5000.000 1391.000    61
+2.19522107E+01+2.48781991E-02-8.44297007E-06+1.30371698E-09-7.53469325E-14    2
-4.34404184E+04-8.34515565E+01+1.20882689E+00+7.78602587E-02-6.16377315E-05    3
+2.60506873E-08-4.52025263E-12-3.66524607E+04+2.64078764E+01+0.00000000E+00    4
BO2C5H10OH 17/8/15      C   5H  11O   3    0G   300.000  5000.000 1395.000    61
+2.28865971E+01+2.40778073E-02-8.16957904E-06+1.26165301E-09-7.29326115E-14    2
-4.48764864E+04-8.92415513E+01+2.71004906E+00+7.28069687E-02-5.37414655E-05    3
+2.08815586E-08-3.34176454E-12-3.80276500E+04+1.85552934E+01+0.00000000E+00    4
CO2C5H10OH 17/8/15      C   5H  11O   3    0G   300.000  5000.000 1406.000    61
+2.22413769E+01+2.43138793E-02-8.17987283E-06+1.25568258E-09-7.22730962E-14    2
-4.13059915E+04-8.36980772E+01-1.39598520E-01+8.39732940E-02-7.03813054E-05    3
+3.10327500E-08-5.52297544E-12-3.42801244E+04+3.38677944E+01+0.00000000E+00    4
IC3H5COCH3 9/ 8/14      C   5H   8O   1    0G   300.000  5000.000 1392.000    31
+1.49935813E+01+1.97788403E-02-6.78313207E-06+1.05481230E-09-6.12614698E-14    2
-2.60877929E+04-5.26202086E+01+1.54292407E+00+5.05432300E-02-3.42434122E-05    3
+1.25252368E-08-1.95302231E-12-2.12702785E+04+1.99855884E+01+0.00000000E+00    4
IC3H5COCH2 9/ 8/14      C   5H   7O   1    0G   300.000  5000.000 1394.000    31
+1.62814836E+01+1.63492954E-02-5.64820836E-06+8.82756224E-10-5.14522209E-14    2
-4.28650692E+03-5.91075528E+01+1.42097745E+00+5.34336638E-02-4.21903633E-05    3
+1.76937615E-08-3.06075290E-12+6.91082980E+02+1.99522060E+01+0.00000000E+00    4
AC3H4COCH3 9/ 8/14      C   5H   7O   1    0G   300.000  5000.000 1384.000    21
+1.60405803E+01+1.62938876E-02-5.49275040E-06+8.45442040E-10-4.87866397E-14    2
-8.30972832E+03-5.83003416E+01+9.48806278E-01+5.17869173E-02-3.74867620E-05    3
+1.40294881E-08-2.14698694E-12-3.10553556E+03+2.26479362E+01+0.00000000E+00    4
NEOC5H12   9/ 8/14      C   5H  12    0    0G   300.000  5000.000 1459.000    41
+2.13410465E+01+2.32500105E-02-8.36387815E-06+1.34306692E-09-7.97752777E-14    2
-3.18056043E+04-1.00649903E+02+8.60482114E-01+4.63444251E-02+2.26557531E-06    3
-1.91739545E-08+6.07291520E-12-2.24020628E+04+1.78235950E+01+0.00000000E+00    4
NEOC5H11   9/ 8/14      C   5H  11    0    0G   300.000  5000.000 1375.000    41
+1.17983312E+01+3.59579648E-02-1.44108662E-05+2.46307665E-09-1.52118262E-13    2
-3.86101387E+03-4.41297337E+01+9.68072098E+00+7.07718151E-03+4.53301778E-05    3
-3.61952123E-08+8.06654396E-12+1.05116941E+03-1.94358274E+01+0.00000000E+00    4
NEOC5H11O2H 9/8/14      C   5H  12O   2    0G   300.000  5000.000 2019.000    61
+2.01975284E+01+2.97380281E-02-1.09930813E-05+1.80338361E-09-1.08851734E-13    2
-3.95165952E+04-8.23753662E+01+3.55225748E-01+6.91131421E-02-3.61242956E-05    3
+6.97537323E-09-9.54855674E-14-3.23388889E+04+2.61109340E+01+0.00000000E+00    4
NEOC5H11O2  9/8/14      C   5H  11O   2    0G   300.000  5000.000 1682.000    51
+1.93713105E+01+2.82612571E-02-1.04670110E-05+1.71917414E-09-1.03854375E-13    2
-2.23544131E+04-7.71662358E+01+1.08144664E+00+6.33534647E-02-3.11938784E-05    3
+4.88883786E-09+2.48584189E-13-1.56455031E+04+2.32475108E+01+0.00000000E+00    4
NEOC5H11O  9/ 8/14      C   5H  11O   1    0G   300.000  5000.000 1374.000    41
+1.47920426E+01+3.60239861E-02-1.44548775E-05+2.47285304E-09-1.52828569E-13    2
-2.12880602E+04-5.86605592E+01+1.11399567E+01+9.95551445E-03+4.37547263E-05    3
-3.60663886E-08+8.13722634E-12-1.57739963E+04-2.54644054E+01+0.00000000E+00    4
NEOC5H10OOH 9/8/14      C   5H  11O   2    0G   300.000  5000.000 1686.000    61
+1.98216577E+01+2.74351153E-02-1.01763800E-05+1.67311287E-09-1.01142157E-13    2
-1.44846637E+04-7.65499851E+01+7.26388728E-01+6.54763558E-02-3.46433563E-05    3
+6.82220142E-09-1.22217205E-13-7.61522056E+03+2.77840799E+01+0.00000000E+00    4
NEO-C5H10O 9/ 8/14      C   5H  10O   1    0G   300.000  5000.000 1465.000    21
+1.88696363E+01+2.18446364E-02-7.48656898E-06+1.16574180E-09-6.78305009E-14    2
-2.76538327E+04-8.33848438E+01-5.80125483E+00+7.19986445E-02-4.12060995E-05    3
+8.52947622E-09+2.15532151E-14-1.85918283E+04+5.13449073E+01+0.00000000E+00    4
NEOC5H10OOH-O2 914      C   5H  11O   4    0G   300.000  5000.000 2038.000    71
+2.43460937E+01+2.84840536E-02-1.05961421E-05+1.74545495E-09-1.05654571E-13    2
-3.35348323E+04-9.58566184E+01+2.12490773E+00+7.51548100E-02-4.39349794E-05    3
+1.09212325E-08-8.06703541E-13-2.57458785E+04+2.47165260E+01+0.00000000E+00    4
NEOC5H9Q2  9/ 8/14      C   5H  11O   4    0G   300.000  5000.000 2050.000    81
+2.48112747E+01+2.76461534E-02-1.03017544E-05+1.69884890E-09-1.02912689E-13    2
-2.56663214E+04-9.64118626E+01+1.90419491E+00+7.68023849E-02-4.67666506E-05    3
+1.25175307E-08-1.11211508E-12-1.77393477E+04+2.75076242E+01+0.00000000E+00    4
NEOC5KET   9/ 8/14      C   5H  10O   3    0G   300.000  5000.000 1396.000    61
+2.11457411E+01+2.34263362E-02-8.03514708E-06+1.24990645E-09-7.26173329E-14    2
-4.99812693E+04-8.04502172E+01+1.99299705E+00+6.63799852E-02-4.41434233E-05    3
+1.47656228E-08-1.97164356E-12-4.31727732E+04+2.30090729E+01+0.00000000E+00    4
NEOC5KETOX 9/ 8/14      C   5H   9O   2    0G   300.000  5000.000 1677.000    41
+1.62834087E+01+2.47667618E-02-8.89982283E-06+1.43325482E-09-8.54232652E-14    2
-2.99100005E+04-5.60198008E+01+3.76958673E+00+4.84037082E-02-2.22215659E-05    3
+2.98251470E-09+2.98064950E-13-2.52993970E+04+1.27918996E+01+0.00000000E+00    4
NEOC5KEJOL 9/ 8/14      C   5H   9O   2    0G   300.000  5000.000 1402.000    51
+1.78858167E+01+2.12423369E-02-7.21947714E-06+1.11609095E-09-6.45625691E-14    2
-3.87680922E+04-6.36233643E+01+1.30298806E+00+5.84132694E-02-3.81961088E-05    3
+1.24622441E-08-1.59437417E-12-3.28976593E+04+2.59154966E+01+0.00000000E+00    4
IC4H6Q2-II 9/ 8/14      C   4H   8O   4    0G   300.000  5000.000 1386.000    61
+2.50360805E+01+1.60230197E-02-5.70704966E-06+9.10412038E-10-5.38294659E-14    2
-2.84196401E+04-9.67186452E+01+2.16408482E-01+8.25572149E-02-7.64540445E-05    3
+3.58211787E-08-6.67718658E-12-2.05694845E+04+3.36943223E+01+0.00000000E+00    4
NEOC5H9O-OOH  9/14      C   5H  10O   3    0G   300.000  5000.000 1429.000    41
+2.34301312E+01+2.26473800E-02-7.84730788E-06+1.22994662E-09-7.18633905E-14    2
-3.86378493E+04-1.00093171E+02-4.33879286E+00+8.23095013E-02-5.24634537E-05    3
+1.40859094E-08-1.00626405E-12-2.87630624E+04+5.04065995E+01+0.00000000E+00    4
C5H10-1                 C   5H  10    0    0G   300.000  5000.000 1390.000    31
+1.43624894E+01+2.26076154E-02-7.70500843E-06+1.19329968E-09-6.91126022E-14    2
-9.99915627E+03-5.12512094E+01-1.65023816E-01+5.30727359E-02-3.10861587E-05    3
+8.92413402E-09-9.81619602E-13-4.57363143E+03+2.80570113E+01+0.00000000E+00    4
C5H10-2    9/ 8/14      C   5H  10    0    0G   300.000  5000.000 1385.000    31
+1.39425521E+01+2.28734997E-02-7.77800113E-06+1.20284861E-09-6.95972140E-14    2
-1.12165700E+04-4.95379542E+01+5.90528835E-01+4.85275113E-02-2.43231598E-05    3
+4.86096027E-09-1.13099201E-13-5.99777644E+03+2.41816377E+01+0.00000000E+00    4
C5H91-1                 C   5H   9    0    0G   300.000  5000.000 1392.000    31
+1.43746526E+01+1.99244772E-02-6.75299634E-06+1.04202761E-09-6.01991076E-14    2
+1.97695686E+04-4.94774744E+01+5.53601698E-01+5.07680916E-02-3.27903964E-05    3
+1.09672330E-08-1.50701628E-12+2.47319519E+04+2.52922332E+01+0.00000000E+00    4
C5H81-3    9/ 8/14      C   5H   8    0    0G   300.000  5000.000 1385.000    21
+1.29945372E+01+1.92678312E-02-6.58966712E-06+1.02295969E-09-5.93441369E-14    2
+4.59040047E+03-4.35689825E+01+1.54882436E+00+4.15042709E-02-2.14359890E-05    3
+4.71145517E-09-2.42142508E-13+9.05636062E+03+1.95665910E+01+0.00000000E+00    4
C5H91-3    9/ 8/14      C   5H   9    0    0G   300.000  5000.000 1390.000    21
+1.39593933E+01+2.09180210E-02-7.14307074E-06+1.10781333E-09-6.42268160E-14    2
+7.02651017E+03-5.03103610E+01-4.68159636E-01+5.13472600E-02-3.05648794E-05    3
+8.82809744E-09-9.61458255E-13+1.23781446E+04+2.83587835E+01+0.00000000E+00    4
C5H91-4    9/ 8/14      C   5H   9    0    0G   300.000  5000.000 1387.000    31
+1.29229725E+01+2.10931621E-02-7.14227112E-06+1.10137556E-09-6.35983966E-14    2
+1.38192408E+04-4.00293126E+01+1.58797615E+00+4.01577239E-02-1.50062687E-05    3
-3.94608061E-10+1.02064182E-12+1.84683983E+04+2.34273438E+01+0.00000000E+00    4
C5H91-5    9/ 8/14      C   5H   9    0    0G   300.000  5000.000 1391.000    31
+1.37334869E+01+2.07003006E-02-7.06962737E-06+1.09638953E-09-6.35591113E-14    2
+1.51176253E+04-4.50794850E+01+2.07676634E-01+4.96049077E-02-3.00621602E-05    3
+9.19962077E-09-1.13246061E-12+2.01251866E+04+2.85856261E+01+0.00000000E+00    4
C5H92-4    9/ 8/14      C   5H   9    0    0G   300.000  5000.000 1384.000    21
+1.35637956E+01+2.11621316E-02-7.20826071E-06+1.11611006E-09-6.46370085E-14    2
+5.82258629E+03-4.87323606E+01+2.55028348E-01+4.69860501E-02-2.40447582E-05    3
+4.89006694E-09-1.15557679E-13+1.09775103E+04+2.46226810E+01+0.00000000E+00    4
C5H92-5    9/ 8/14      C   5H   9    0    0G   300.000  5000.000 1386.000    31
+1.32988753E+01+2.09845923E-02-7.14999241E-06+1.10717347E-09-6.41183619E-14    2
+1.39270369E+04-4.32758927E+01+9.96363945E-01+4.49148898E-02-2.30951498E-05    3
+5.01698735E-09-2.38646470E-13+1.87161506E+04+2.45616052E+01+0.00000000E+00    4
C5H9O1-3   9/ 8/14      C   5H   9O   1    0G   300.000  5000.000 1379.000    31
+1.78860333E+01+2.04837367E-02-7.16613461E-06+1.12948597E-09-6.62221468E-14    2
-4.33139568E+03-6.72851315E+01+2.49666166E+00+5.20326105E-02-3.09828268E-05    3
+9.02567482E-09-1.04311127E-12+1.54758549E+03+1.70868328E+01+0.00000000E+00    4
C5H9O2-4   9/ 8/14      C   5H   9O   1    0G   300.000  5000.000 1376.000    31
+1.73707371E+01+2.09044827E-02-7.30723872E-06+1.15106814E-09-6.74601377E-14    2
-5.48020434E+03-6.50109045E+01+3.38899911E+00+4.71704753E-02-2.40389823E-05    3
+4.99166621E-09-2.03242522E-13+1.15232772E+02+1.25183625E+01+0.00000000E+00    4
BC5H10     9/ 8/14      C   5H  10    0    0G   300.000  5000.000 1389.000    31
+1.40426423E+01+2.27915348E-02-7.74902598E-06+1.19814522E-09-6.93127003E-14    2
-1.32160483E+04-5.14469569E+01+6.04882839E-01+4.96635256E-02-2.66571142E-05    3
+6.47312078E-09-4.84017883E-13-8.06312207E+03+2.23818263E+01+0.00000000E+00    4
CC5H10     9/ 8/14      C   5H  10    0    0G   300.000  5000.000 1394.000    31
+1.44242929E+01+2.26454984E-02-7.73646334E-06+1.19999861E-09-6.95711276E-14    2
-1.14981027E+04-5.30391197E+01-9.64397004E-01+5.68482691E-02-3.66324275E-05    3
+1.23008921E-08-1.71392531E-12-5.93502026E+03+3.02998433E+01+0.00000000E+00    4
CC5H9-A                 C   5H   9    0    0G   300.000  5000.000 1393.000    31
+1.38635892E+01+2.06362872E-02-7.05717373E-06+1.09539676E-09-6.35381849E-14    2
+1.36104251E+04-4.72507189E+01-6.78909715E-01+5.37496002E-02-3.61116825E-05    3
+1.28563411E-08-1.92155723E-12+1.87974429E+04+3.12403382E+01+0.00000000E+00    4
CC5H9-B    9/ 8/14      C   5H   9    0    0G   300.000  5000.000 1392.000    21
+1.35249511E+01+2.14363755E-02-7.35304116E-06+1.14368637E-09-6.64363518E-14    2
+5.41381916E+03-5.00302394E+01-6.91501860E-01+5.09804846E-02-2.96448293E-05    3
+8.28273022E-09-8.57575066E-13+1.07478467E+04+2.76711552E+01+0.00000000E+00    4
AC5H9O-C                C   5H   9O   1    0G   300.000  5000.000 1382.000    31
+1.76789601E+01+2.05915073E-02-7.18764438E-06+1.13116483E-09-6.62505034E-14    2
-6.25146818E+03-6.62131721E+01+2.04951318E+00+5.36584877E-02-3.35086710E-05    3
+1.06174235E-08-1.39224338E-12-3.85112518E+02+1.91077262E+01+0.00000000E+00    4
CC5H9O-B   9/ 8/14      C   5H   9O   1    0G   300.000  5000.000 1377.000    31
+1.86974377E+01+1.84542537E-02-6.18682537E-06+9.48850967E-10-5.46203980E-14    2
-7.15897769E+03-7.26540429E+01+2.75614808E+00+5.20514036E-02-3.10966938E-05    3
+8.25895065E-09-6.59917121E-13-1.35162741E+03+1.40990119E+01+0.00000000E+00    4
AC5H10                  C   5H  10    0    0G   300.000  5000.000 1392.000    31
+1.41931279E+01+2.26551019E-02-7.70008627E-06+1.19031326E-09-6.88489604E-14    2
-1.19491010E+04-5.10688681E+01-5.39429136E-01+5.44489715E-02-3.32707895E-05    3
+1.03047694E-08-1.28363329E-12-6.53967251E+03+2.90349986E+01+0.00000000E+00    4
AC5H9-A2                C   5H   9    0    0G   300.000  5000.000 1385.000    21
+1.50019889E+01+1.95965428E-02-6.60205927E-06+1.01535593E-09-5.85454957E-14    2
+5.90081014E+03-5.54528992E+01-9.54047710E-01+5.50153471E-02-3.58307910E-05    3
+1.16444141E-08-1.49086833E-12+1.15959514E+04+3.08476806E+01+0.00000000E+00    4
AC5H9-C                 C   5H   9    0    0G   300.000  5000.000 1392.000    21
+1.37918110E+01+2.09644966E-02-7.13793293E-06+1.10480881E-09-6.39628018E-14    2
+5.09555600E+03-5.01391436E+01-8.41372657E-01+5.27157283E-02-3.27334707E-05    3
+1.01974035E-08-1.26084730E-12+1.04321036E+04+2.93316754E+01+0.00000000E+00    4
AC5H9-D                 C   5H   9    0    0G   300.000  5000.000 1393.000    31
+1.35607521E+01+2.07514878E-02-7.06608626E-06+1.09362345E-09-6.33083050E-14    2
+1.31896844E+04-4.48718988E+01-1.67398152E-01+5.09876974E-02-3.22615638E-05    3
+1.05911843E-08-1.43705463E-12+1.81792947E+04+2.95710715E+01+0.00000000E+00    4
B2E2M1OJ                C   5H   9O   1    0G   300.000  5000.000 2003.000    31
+1.35666458E+01+2.56547934E-02-9.37226256E-06+1.52518398E-09-9.15378763E-14    2
-3.58767067E+03-4.27272791E+01+5.64762692E+00+3.43609862E-02-5.60649548E-06    3
-5.19111402E-09+1.73155461E-12-6.65737793E+00+3.13825267E+00+0.00000000E+00    4
B13DE2M                 C   5H   8    0    0G   300.000  5000.000 1397.000    21
+1.40757545E+01+1.82375566E-02-6.20747687E-06+9.60350919E-10-5.55741525E-14    2
+2.40033881E+03-5.12988284E+01-4.72170009E-01+5.59413257E-02-4.50458826E-05    3
+1.96181377E-08-3.52009647E-12+7.14960489E+03+2.56276807E+01+0.00000000E+00    4
B13DE2MJ                C   5H   7    0    0G   300.000  5000.000 1393.000    11
+1.48413344E+01+1.52425753E-02-5.13559858E-06+7.89787260E-10-4.55353492E-14    2
+2.02661570E+04-5.54474955E+01-8.98037227E-01+5.65174321E-02-4.76107829E-05    3
+2.09672106E-08-3.73076319E-12+2.52881763E+04+2.74966602E+01+0.00000000E+00    4
B12DE3M   11/12/12 THERMC   5H   8    0    0G   300.000  5000.000 1388.000    21
+1.37093177E+01+1.85726726E-02-6.33115904E-06+9.80719059E-10-5.68099894E-14    2
+8.59518752E+03-4.88749621E+01+1.27860173E+00+4.54917474E-02-2.82334169E-05    3
+8.98449372E-09-1.17220042E-12+1.31637341E+04+1.87039373E+01+0.00000000E+00    4
B2E3M1OJ                C   5H   9O   1    0G   300.000  5000.000 2003.000    31
+1.35666458E+01+2.56547934E-02-9.37226256E-06+1.52518398E-09-9.15378763E-14    2
-3.58767067E+03-4.27272791E+01+5.64762692E+00+3.43609862E-02-5.60649548E-06    3
-5.19111402E-09+1.73155461E-12-6.65737793E+00+3.13825267E+00+0.00000000E+00    4
TC4H8CHO   9/ 7/95 THERMC   5H   9O   1    0G   300.000  5000.000 1397.00     41
+1.79663933E+01+1.94207117E-02-6.67409451E-06+1.03969221E-09-6.04702651E-14    2
-1.33368585E+04-6.79819424E+01-9.58078294E-01+6.42003258E-02-4.70776827E-05    3
+1.75737698E-08-2.64896151E-12-6.86582501E+03+3.33781112E+01+0.00000000E+00    4
O2C4H8CHO  9/ 7/95 THERMC   5H   9O   3    0G   300.000  5000.000 1395.00     51
+2.12629904E+01+2.14072282E-02-7.38342949E-06+1.15281523E-09-6.71508438E-14    2
-3.16854524E+04-7.99828703E+01+1.91847699E+00+6.67245869E-02-4.80871046E-05    3
+1.78588690E-08-2.71163880E-12-2.49837984E+04+2.38577867E+01+0.00000000E+00    4
O2HC4H8CO  9/ 7/95 THERMC   5H   9O   3    0G   300.000  5000.000 1394.00     61
+2.38219630E+01+1.91411448E-02-6.67919154E-06+1.05127303E-09-6.15876805E-14    2
-3.23093973E+04-9.42580755E+01+1.82607262E+00+6.93466111E-02-4.93125140E-05    3
+1.69848340E-08-2.26117657E-12-2.46578311E+04+2.41167544E+01+0.00000000E+00    4
PC4H9CHO                C   5H  10O   1    0G   300.000  5000.000 1383.000    41
+1.71928366E+01+2.24205079E-02-7.66524563E-06+1.18999819E-09-6.90481012E-14    2
-3.62048450E+04-6.39265450E+01+1.55168051E+00+5.17580624E-02-2.47521866E-05    3
+3.39585733E-09+4.54214964E-13-3.01104924E+04+2.25340321E+01+0.00000000E+00    4
PC4H9CO                 C   5H   9O   1    0G   300.000  5000.000 1380.000    41
+1.67761337E+01+2.02898448E-02-6.94418179E-06+1.07888297E-09-6.26360391E-14    2
-1.72426942E+04-6.00185187E+01+2.32674439E+00+4.69567990E-02-2.17002843E-05    3
+2.33166983E-09+6.15109331E-13-1.15824032E+04+1.99866279E+01+0.00000000E+00    4
PC4H8CHO-1              C   5H   9O   1    0G   300.000  5000.000 1391.000    41
+1.73203841E+01+2.00050584E-02-6.88462599E-06+1.07357298E-09-6.24869113E-14    2
-1.60879440E+04-6.51443168E+01+8.84469923E-01+5.26232725E-02-2.83373818E-05    3
+5.66303879E-09-3.63459101E-15-9.89241254E+03+2.50250388E+01+0.00000000E+00    4
PC4H8CHO-2              C   5H   9O   1    0G   300.000  5000.000 1426.000    41
+1.58456286E+01+2.08430527E-02-7.08562851E-06+1.09605491E-09-6.34445999E-14    2
-1.24300179E+04-5.32908403E+01+3.19129086E+00+3.91487154E-02-8.88573585E-06    3
-5.86340400E-09+2.44961462E-12-7.02633915E+03+1.84682536E+01+0.00000000E+00    4
PC4H8CHO-3              C   5H   9O   1    0G   300.000  5000.000 1426.000    41
+1.58456286E+01+2.08430527E-02-7.08562851E-06+1.09605491E-09-6.34445999E-14    2
-1.24300179E+04-5.32908403E+01+3.19129086E+00+3.91487154E-02-8.88573585E-06    3
-5.86340400E-09+2.44961462E-12-7.02633915E+03+1.84682536E+01+0.00000000E+00    4
PC4H8CHO-4              C   5H   9O   1    0G   300.000  5000.000 1383.000    41
+1.66333143E+01+2.03619734E-02-6.95844731E-06+1.08002411E-09-6.26591600E-14    2
-1.10824930E+04-5.81167187E+01+1.89962807E+00+4.83598549E-02-2.37381500E-05    3
+3.58762168E-09+3.40201608E-13-5.38702187E+03+2.31840311E+01+0.00000000E+00    4
AC3H5CHO                C   4H   6O   1    0G   300.000  5000.000 1387.000    21
+1.27609075E+01+1.48416812E-02-5.16797249E-06+8.12052956E-10-4.75111888E-14    2
-1.54802190E+04-4.05362549E+01-1.35627837E-01+4.32102800E-02-2.86018998E-05    3
+9.48372797E-09-1.26553781E-12-1.08101418E+04+2.93765145E+01+0.00000000E+00    4
PC4H8CHO-1O2 10/8/15    C   5H   9O   3    0G   300.000  5000.000 1385.000    51
+2.46719452E+01+1.85504127E-02-6.42209840E-06+1.00647312E-09-5.88171032E-14    2
-3.18555321E+04-9.71440808E+01-4.63291072E-01+8.02504798E-02-6.47236563E-05    3
+2.62037194E-08-4.25127975E-12-2.34955268E+04+3.66761324E+01+0.00000000E+00    4
PC4H8CHO-2O2 10/8/15    C   5H   9O   3    0G   300.000  5000.000 1404.000    51
+2.16725120E+01+2.03883823E-02-6.89025420E-06+1.06159257E-09-6.12789415E-14    2
-3.20581874E+04-8.08233009E+01+3.75698588E+00+5.99220385E-02-3.84711370E-05    3
+1.16653123E-08-1.26664695E-12-2.57207120E+04+1.60217605E+01+0.00000000E+00    4
PC4H8CHO-3O2 10/8/15    C   5H   9O   3    0G   300.000  5000.000 1404.000    51
+2.16725120E+01+2.03883823E-02-6.89025420E-06+1.06159257E-09-6.12789415E-14    2
-3.20581874E+04-8.08233009E+01+3.75698588E+00+5.99220385E-02-3.84711370E-05    3
+1.16653123E-08-1.26664695E-12-2.57207120E+04+1.60217605E+01+0.00000000E+00    4
PC4H8CHO-4O2 10/8/15    C   5H   9O   3    0G   300.000  5000.000 1385.000    51
+2.12856144E+01+2.12771293E-02-7.31814716E-06+1.14082494E-09-6.63900040E-14    2
-3.02079416E+04-7.82029614E+01+3.37850952E+00+5.77659231E-02-3.28975023E-05    3
+7.80995858E-09-4.14571925E-13-2.35309122E+04+1.97380195E+01+0.00000000E+00    4
C4H7CHO-2  10/8/15 THERMC   5H   8O   1    0G   300.000  5000.000 1390.000    31
+1.62588601E+01+1.87787531E-02-6.45805165E-06+1.00641261E-09-5.85466414E-14    2
-2.44023233E+04-5.96450353E+01+3.69688874E-04+5.71382743E-02-4.15287925E-05    3
+1.58289787E-08-2.49867087E-12-1.87655817E+04+2.75869712E+01+0.00000000E+00    4
C4H7CHO-2               C   5H   8O   1    0G   300.000  5000.000 1390.000    31
+1.62588601E+01+1.87787531E-02-6.45805165E-06+1.00641261E-09-5.85466414E-14    2
-2.44023233E+04-5.96450353E+01+3.69688874E-04+5.71382743E-02-4.15287925E-05    3
+1.58289787E-08-2.49867087E-12-1.87655817E+04+2.75869712E+01+0.00000000E+00    4
C4H7CHO-2  10/8/15 THERMC   5H   8O   1    0G   300.000  5000.000 1390.000    31
+1.62588601E+01+1.87787531E-02-6.45805165E-06+1.00641261E-09-5.85466414E-14    2
-2.44023233E+04-5.96450353E+01+3.69688874E-04+5.71382743E-02-4.15287925E-05    3
+1.58289787E-08-2.49867087E-12-1.87655817E+04+2.75869712E+01+0.00000000E+00    4
C4H7CHO-2               C   5H   8O   1    0G   300.000  5000.000 1390.000    31
+1.62588601E+01+1.87787531E-02-6.45805165E-06+1.00641261E-09-5.85466414E-14    2
-2.44023233E+04-5.96450353E+01+3.69688874E-04+5.71382743E-02-4.15287925E-05    3
+1.58289787E-08-2.49867087E-12-1.87655817E+04+2.75869712E+01+0.00000000E+00    4
C4H7CHO-2  10/8/15 THERMC   5H   8O   1    0G   300.000  5000.000 1390.000    31
+1.62588601E+01+1.87787531E-02-6.45805165E-06+1.00641261E-09-5.85466414E-14    2
-2.44023233E+04-5.96450353E+01+3.69688874E-04+5.71382743E-02-4.15287925E-05    3
+1.58289787E-08-2.49867087E-12-1.87655817E+04+2.75869712E+01+0.00000000E+00    4
C4H7CHO-2               C   5H   8O   1    0G   300.000  5000.000 1390.000    31
+1.62588601E+01+1.87787531E-02-6.45805165E-06+1.00641261E-09-5.85466414E-14    2
-2.44023233E+04-5.96450353E+01+3.69688874E-04+5.71382743E-02-4.15287925E-05    3
+1.58289787E-08-2.49867087E-12-1.87655817E+04+2.75869712E+01+0.00000000E+00    4
C4H7CHO-2  10/8/15 THERMC   5H   8O   1    0G   300.000  5000.000 1390.000    31
+1.62588601E+01+1.87787531E-02-6.45805165E-06+1.00641261E-09-5.85466414E-14    2
-2.44023233E+04-5.96450353E+01+3.69688874E-04+5.71382743E-02-4.15287925E-05    3
+1.58289787E-08-2.49867087E-12-1.87655817E+04+2.75869712E+01+0.00000000E+00    4
C4H7CHO-2               C   5H   8O   1    0G   300.000  5000.000 1390.000    31
+1.62588601E+01+1.87787531E-02-6.45805165E-06+1.00641261E-09-5.85466414E-14    2
-2.44023233E+04-5.96450353E+01+3.69688874E-04+5.71382743E-02-4.15287925E-05    3
+1.58289787E-08-2.49867087E-12-1.87655817E+04+2.75869712E+01+0.00000000E+00    4
C4H7CHO-2  10/8/15 THERMC   5H   8O   1    0G   300.000  5000.000 1390.000    31
+1.62588601E+01+1.87787531E-02-6.45805165E-06+1.00641261E-09-5.85466414E-14    2
-2.44023233E+04-5.96450353E+01+3.69688874E-04+5.71382743E-02-4.15287925E-05    3
+1.58289787E-08-2.49867087E-12-1.87655817E+04+2.75869712E+01+0.00000000E+00    4
C4H7CHO-2               C   5H   8O   1    0G   300.000  5000.000 1390.000    31
+1.62588601E+01+1.87787531E-02-6.45805165E-06+1.00641261E-09-5.85466414E-14    2
-2.44023233E+04-5.96450353E+01+3.69688874E-04+5.71382743E-02-4.15287925E-05    3
+1.58289787E-08-2.49867087E-12-1.87655817E+04+2.75869712E+01+0.00000000E+00    4
C4H7CHO-2  10/8/15 THERMC   5H   8O   1    0G   300.000  5000.000 1390.000    31
+1.62588601E+01+1.87787531E-02-6.45805165E-06+1.00641261E-09-5.85466414E-14    2
-2.44023233E+04-5.96450353E+01+3.69688874E-04+5.71382743E-02-4.15287925E-05    3
+1.58289787E-08-2.49867087E-12-1.87655817E+04+2.75869712E+01+0.00000000E+00    4
C4H7CHO-2               C   5H   8O   1    0G   300.000  5000.000 1390.000    31
+1.62588601E+01+1.87787531E-02-6.45805165E-06+1.00641261E-09-5.85466414E-14    2
-2.44023233E+04-5.96450353E+01+3.69688874E-04+5.71382743E-02-4.15287925E-05    3
+1.58289787E-08-2.49867087E-12-1.87655817E+04+2.75869712E+01+0.00000000E+00    4
C4H7CHO-2  10/8/15 THERMC   5H   8O   1    0G   300.000  5000.000 1390.000    31
+1.62588601E+01+1.87787531E-02-6.45805165E-06+1.00641261E-09-5.85466414E-14    2
-2.44023233E+04-5.96450353E+01+3.69688874E-04+5.71382743E-02-4.15287925E-05    3
+1.58289787E-08-2.49867087E-12-1.87655817E+04+2.75869712E+01+0.00000000E+00    4
C4H7CHO-2               C   5H   8O   1    0G   300.000  5000.000 1390.000    31
+1.62588601E+01+1.87787531E-02-6.45805165E-06+1.00641261E-09-5.85466414E-14    2
-2.44023233E+04-5.96450353E+01+3.69688874E-04+5.71382743E-02-4.15287925E-05    3
+1.58289787E-08-2.49867087E-12-1.87655817E+04+2.75869712E+01+0.00000000E+00    4
C4H7CHO-2  10/8/15 THERMC   5H   8O   1    0G   300.000  5000.000 1390.000    31
+1.62588601E+01+1.87787531E-02-6.45805165E-06+1.00641261E-09-5.85466414E-14    2
-2.44023233E+04-5.96450353E+01+3.69688874E-04+5.71382743E-02-4.15287925E-05    3
+1.58289787E-08-2.49867087E-12-1.87655817E+04+2.75869712E+01+0.00000000E+00    4
C4H7CHO-2               C   5H   8O   1    0G   300.000  5000.000 1390.000    31
+1.62588601E+01+1.87787531E-02-6.45805165E-06+1.00641261E-09-5.85466414E-14    2
-2.44023233E+04-5.96450353E+01+3.69688874E-04+5.71382743E-02-4.15287925E-05    3
+1.58289787E-08-2.49867087E-12-1.87655817E+04+2.75869712E+01+0.00000000E+00    4
C4H7CHO-3  10/8/15 THERMC   5H   8O   1    0G   300.000  5000.000 1385.000    31
+1.55930799E+01+1.96344789E-02-6.81722246E-06+1.06912344E-09-6.24665079E-14    2
-2.08408048E+04-5.47830431E+01+4.14190085E-01+5.12150376E-02-3.06682310E-05    3
+8.72168876E-09-9.15725235E-13-1.51552520E+04+2.81574532E+01+0.00000000E+00    4
C4H7CHO-4  10/8/15 THERMC   5H   8O   1    0G   300.000  5000.000 2020.000    31
+1.37156197E+01+2.16425024E-02-7.67112142E-06+1.22483309E-09-7.25906717E-14    2
-1.91110565E+04-4.33806662E+01+1.15814338E+00+4.81746752E-02-2.67363172E-05    3
+6.50396537E-09-4.78416928E-13-1.47390215E+04+2.46792248E+01+0.00000000E+00    4
NC3H7COCH3 10/6/15 THERMC   5H  10O   1    0G   300.000  5000.000 1387.000    41
+1.59632618E+01+2.26394805E-02-7.56430418E-06+1.15632032E-09-6.63757297E-14    2
-3.92822369E+04-5.65033421E+01+2.22465879E+00+4.82791863E-02-2.21019858E-05    3
+2.64029906E-09+5.23720489E-13-3.39379060E+04+1.94495002E+01+0.00000000E+00    4
C2H5COC2H5 10/6/15 THERMC   5H  10O   1    0G   300.000  5000.000 1421.000    41
+1.65155931E+01+2.18966306E-02-7.26184066E-06+1.10537530E-09-6.32910022E-14    2
-3.96722497E+04-6.11243728E+01+3.04335984E+00+4.24811577E-02-1.12087588E-05    3
-5.05051822E-09+2.35367193E-12-3.40615638E+04+1.48305047E+01+0.00000000E+00    4
NC3H7COCH2 10/6/15 THERMC   5H   9O   1    0G   300.000  5000.000 1393.000    41
+1.72611127E+01+1.91828746E-02-6.41680319E-06+9.82027213E-10-5.64270287E-14    2
-1.74829806E+04-6.30397964E+01+2.14964962E+00+5.09715972E-02-2.97744827E-05    3
+7.64275255E-09-5.47753503E-13-1.19838512E+04+1.91969246E+01+0.00000000E+00    4
CH3CH2CHCOCH3 10/6/15   C   5H   9O   1    0G   300.000  5000.000 1428.000    41
+1.53040392E+01+2.03924168E-02-6.74389287E-06+1.02444156E-09-5.85693457E-14    2
-1.95765010E+04-4.96835091E+01+3.62180151E+00+3.78869197E-02-9.52099354E-06    3
-4.70140858E-09+2.11456934E-12-1.46643385E+04+1.63246571E+01+0.00000000E+00    4
CH3CHCH2COCH3 10/6/15   C   5H   9O   1    0G   300.000  5000.000 1313.000    41
+1.45647685E+01+2.10276788E-02-6.95711397E-06+1.05654321E-09-6.03737583E-14    2
-1.54618001E+04-4.55117654E+01+3.82775077E+00+3.59153332E-02-6.78571299E-06    3
-6.24819689E-09+2.43917244E-12-1.08496104E+04+1.55399306E+01+0.00000000E+00    4
CH2CH2CH2COCH3 10/6/15  C   5H   9O   1    0G   300.000  5000.000 2010.000    41
+1.36121876E+01+2.29083157E-02-7.89568575E-06+1.23743112E-09-7.24018569E-14    2
-1.31339181E+04-4.00994585E+01+2.03928898E+00+4.76715898E-02-2.60373643E-05    3
+6.44110554E-09-5.11322699E-13-9.14243040E+03+2.25010591E+01+0.00000000E+00    4
CH2CH2COC2H5 10/6/15    C   5H   9O   1    0G   300.000  5000.000 1418.000    41
+1.58030158E+01+2.00450814E-02-6.64102020E-06+1.01015297E-09-5.78091691E-14    2
-1.44839773E+04-5.37408145E+01+3.36988365E+00+3.93333507E-02-1.08692381E-05    3
-4.28049004E-09+2.08635748E-12-9.33794632E+03+1.62475992E+01+0.00000000E+00    4
CH3CHCOC2H5 10/6/15     C   5H   9O   1    0G   300.000  5000.000 1426.000    41
+1.52590939E+01+2.06874083E-02-6.90185396E-06+1.05491074E-09-6.05775562E-14    2
-1.97701234E+04-5.03404450E+01+4.26150430E+00+3.32446421E-02-1.19632509E-06    3
-1.01813061E-08+3.34232716E-12-1.47673892E+04+1.31662371E+01+0.00000000E+00    4
NC52ONEO2-3 10/8/15     C   5H   9O   3    0G   300.000  5000.000 1389.000    51
+2.32384890E+01+1.91383699E-02-6.48795686E-06+1.00265179E-09-5.80286197E-14    2
-3.48643643E+04-8.86014914E+01+3.67212944E-01+7.61782682E-02-6.13904833E-05    3
+2.51922695E-08-4.15673555E-12-2.73490750E+04+3.28428407E+01+0.00000000E+00    4
NC52ONEO2-4 10/8/15     C   5H   9O   3    0G   300.000  5000.000 1419.000    51
+2.05185681E+01+2.04863743E-02-6.73858014E-06+1.01931995E-09-5.80865415E-14    2
-3.51672453E+04-7.38258122E+01+4.46745059E+00+5.62677767E-02-3.55388942E-05    3
+1.07130185E-08-1.15039744E-12-2.95536320E+04+1.27650471E+01+0.00000000E+00    4
NC52ONEO2-5 10/8/15     C   5H   9O   3    0G   300.000  5000.000 1388.000    51
+2.00576970E+01+2.15456046E-02-7.24499615E-06+1.11255956E-09-6.40750213E-14    2
-3.33006712E+04-7.08203167E+01+4.08984713E+00+5.40452788E-02-2.97970958E-05    3
+6.76825508E-09-2.84375003E-13-2.73624576E+04+1.64944454E+01+0.00000000E+00    4
NC53ONEO2-1 10/8/15     C   5H   9O   3    0G   300.000  5000.000 1472.000    51
+2.08297563E+01+2.14528808E-02-7.34744816E-06+1.14331164E-09-6.64861408E-14    2
-3.41829302E+04-7.69526850E+01+4.51723400E+00+4.63561824E-02-1.26143575E-05    3
-5.62683827E-09+2.63012314E-12-2.73321757E+04+1.51181731E+01+0.00000000E+00    4
NC53ONEO2-2 10/8/15     C   5H   9O   3    0G   300.000  5000.000 1386.000    51
+2.33146573E+01+1.91100357E-02-6.48744531E-06+1.00363367E-09-5.81318155E-14    2
-3.50527575E+04-8.98266438E+01+1.18594239E+00+7.06410637E-02-5.13727958E-05    3
+1.83400895E-08-2.55856018E-12-2.74781465E+04+2.88673640E+01+0.00000000E+00    4
NC52ONE-3 10/ 8/15 THERMC   5H   8O   1    0G   300.000  5000.000 1388.000    31
+1.48312595E+01+2.01259287E-02-6.94970483E-06+1.08573546E-09-6.32625551E-14    2
-2.65938915E+04-5.14361841E+01+8.18407003E-01+5.17195551E-02-3.47852250E-05    3
+1.26179448E-08-1.96289033E-12-2.15095891E+04+2.44001463E+01+0.00000000E+00    4
NC52ONE-4 10/ 8/15 THERMC   5H   8O   1    0G   300.000  5000.000 1395.000    31
+1.45047399E+01+1.99954720E-02-6.81519480E-06+1.05547414E-09-6.11274397E-14    2
-2.26071842E+04-4.74948237E+01+2.46588134E-01+5.27913864E-02-3.58755256E-05    3
+1.29117478E-08-1.94285390E-12-1.75679347E+04+2.93219925E+01+0.00000000E+00    4
NC53ONE-1 10/ 8/15 THERMC   5H   8O   1    0G   300.000  5000.000 1388.000    31
+1.54699471E+01+1.94419026E-02-6.68487150E-06+1.04158457E-09-6.05841804E-14    2
-2.56037925E+04-5.50815753E+01+1.06845510E+00+4.97050279E-02-2.97718118E-05    3
+8.51066096E-09-8.95411427E-13-2.02580056E+04+2.34730078E+01+0.00000000E+00    4
NC5H11OH  10/ 7/15 THERMC   5H  12O   1    0G   300.000  5000.000 1399.000    51
+1.81326422E+01+2.58734469E-02-8.76147510E-06+1.35108218E-09-7.80169568E-14    2
-4.49393846E+04-6.77258765E+01-7.40082992E-01+6.83880275E-02-4.47177434E-05    3
+1.49115071E-08-1.99981896E-12-3.82501077E+04+3.41515985E+01+0.00000000E+00    4
C5H10OH11 10/ 7/15 THERMC   5H  11O   1    0G   300.000  5000.000 1394.000    51
+1.80953018E+01+2.33361161E-02-7.88463541E-06+1.21428332E-09-7.00616136E-14    2
-2.30206675E+04-6.61675776E+01+4.26049537E-01+6.31258286E-02-4.15122762E-05    3
+1.38895665E-08-1.86732010E-12-1.67596661E+04+2.92144309E+01+0.00000000E+00    4
C5H10OH12 10/ 7/15 THERMC   5H  11O   1    0G   300.000  5000.000 1394.000    51
+1.71780951E+01+2.42601001E-02-8.22986526E-06+1.27049816E-09-7.34155598E-14    2
-2.04290445E+04-5.93472290E+01+1.84753679E+00+5.73086840E-02-3.47271444E-05    3
+1.06516140E-08-1.30777652E-12-1.47995754E+04+2.40150308E+01+0.00000000E+00    4
C5H10OH13 10/ 7/15 THERMC   5H  11O   1    0G   300.000  5000.000 1402.000    51
+1.68143234E+01+2.44876194E-02-8.29372543E-06+1.27921101E-09-7.38804613E-14    2
-2.12567818E+04-5.74573295E+01+5.41167710E-01+5.66862244E-02-2.94678472E-05    3
+5.84904634E-09-3.31866473E-14-1.50943752E+04+3.18827466E+01+0.00000000E+00    4
C5H10OH14 10/ 7/15 THERMC   5H  11O   1    0G   300.000  5000.000 1402.000    51
+1.68143234E+01+2.44876194E-02-8.29372543E-06+1.27921101E-09-7.38804613E-14    2
-2.12567818E+04-5.74573295E+01+5.41167710E-01+5.66862244E-02-2.94678472E-05    3
+5.84904634E-09-3.31866473E-14-1.50943752E+04+3.18827466E+01+0.00000000E+00    4
C5H10OH15 10/ 7/15 THERMC   5H  11O   1    0G   300.000  5000.000 1400.000    51
+1.74868543E+01+2.39842944E-02-8.13298324E-06+1.25529418E-09-7.25301446E-14    2
-1.97969015E+04-6.14612340E+01-3.94307021E-01+6.50012333E-02-4.38043364E-05    3
+1.52539819E-08-2.16516288E-12-1.35258816E+04+3.48138101E+01+0.00000000E+00    4
C5H10OH-1O2    10/ 8/15 C   5H  11O   3    0G   300.000  5000.000 1396.000    61
+2.29458771E+01+2.45179524E-02-8.42764796E-06+1.31282727E-09-7.63477543E-14    2
-4.34982351E+04-8.92569973E+01+1.87266560E+00+7.35120790E-02-5.19769726E-05    3
+1.89528387E-08-2.82611232E-12-3.61605500E+04+2.39948500E+01+0.00000000E+00    4
C5H10OH-2O2    10/ 8/15 C   5H  11O   3    0G   300.000  5000.000 1406.000    61
+2.28162462E+01+2.40750309E-02-8.15387271E-06+1.25759554E-09-7.26292545E-14    2
-4.09893865E+04-8.60865796E+01+1.54218231E+00+7.57844091E-02-5.63028041E-05    3
+2.16374600E-08-3.37143496E-12-3.38651232E+04+2.73478003E+01+0.00000000E+00    4
C5H10OH-3O2    10/ 8/15 C   5H  11O   3    0G   300.000  5000.000 1406.000    61
+2.28162462E+01+2.40750309E-02-8.15387271E-06+1.25759554E-09-7.26292545E-14    2
-4.09893865E+04-8.60865796E+01+1.54218231E+00+7.57844091E-02-5.63028041E-05    3
+2.16374600E-08-3.37143496E-12-3.38651232E+04+2.73478003E+01+0.00000000E+00    4
C5H10OH-4O2    10/ 8/15 C   5H  11O   3    0G   300.000  5000.000 1406.000    61
+2.28162462E+01+2.40750309E-02-8.15387271E-06+1.25759554E-09-7.26292545E-14    2
-4.09893865E+04-8.60865796E+01+1.54218231E+00+7.57844091E-02-5.63028041E-05    3
+2.16374600E-08-3.37143496E-12-3.38651232E+04+2.73478003E+01+0.00000000E+00    4
C5H10OH-5O2    10/ 8/15 C   5H  11O   3    0G   300.000  5000.000 1397.000    61
+2.21449702E+01+2.49621926E-02-8.52928879E-06+1.32336610E-09-7.67473293E-14    2
-3.89467600E+04-8.16310639E+01+1.13788816E+00+7.41287041E-02-5.25165329E-05    3
+1.92381362E-08-2.87963457E-12-3.16767835E+04+3.11292521E+01+0.00000000E+00    4
C5H9OH1-1     10/ 8/15  C   5H  10O   1    0G   300.000  5000.000 1401.000    41
+1.75799784E+01+2.15510873E-02-7.24423039E-06+1.11154167E-09-6.39602647E-14    2
-3.19843372E+04-6.59853552E+01-7.52968139E-01+6.84304063E-02-5.40649298E-05    3
+2.26640783E-08-3.88274568E-12-2.60259987E+04+3.10300945E+01+0.00000000E+00    4
C5H9OH1-2     10/ 8/15  C   5H  10O   1    0G   300.000  5000.000 1375.000    41
+1.62865282E+01+2.40392163E-02-8.40885938E-06+1.32515728E-09-7.76837502E-14    2
-2.99434873E+04-5.80985901E+01+1.71304900E+00+5.05617859E-02-2.46539338E-05    3
+4.87081503E-09-1.89220960E-13-2.39589376E+04+2.31277850E+01+0.00000000E+00    4
C5H9OH1-3     10/ 8/15  C   5H  10O   1    0G   300.000  5000.000 1391.000    41
+1.62749224E+01+2.27984390E-02-7.70751766E-06+1.18747528E-09-6.85336287E-14    2
-3.02380128E+04-5.75828357E+01+1.88732713E-01+5.71777712E-02-3.44214841E-05    3
+9.99837019E-09-1.07315871E-12-2.43560647E+04+2.99036243E+01+0.00000000E+00    4
C5H9OH1-4     10/ 8/15  C   5H  10O   1    0G   300.000  5000.000 1396.000    41
+1.66790471E+01+2.25496587E-02-7.64069183E-06+1.17887585E-09-6.81025445E-14    2
-2.90316501E+04-5.92057123E+01-5.42247537E-01+6.16234351E-02-4.10470356E-05    3
+1.39787947E-08-1.92326047E-12-2.29560111E+04+3.36582311E+01+0.00000000E+00    4
NC6H14                  C   6H  14    0    0G   300.000  5000.000 1394.000    51
+1.91649837E+01+3.02733796E-02-1.03172746E-05+1.59774518E-09-9.25291178E-14    2
-3.01230801E+04-7.69633109E+01-6.06787842E-01+7.23956364E-02-4.33845424E-05    3
+1.28945357E-08-1.49361322E-12-2.28192378E+04+3.07154747E+01+0.00000000E+00    4
C6H13-1                 C   6H  13    0    0G   300.000  5000.000 1395.000    51
+1.85287088E+01+2.83718554E-02-9.68391797E-06+1.50116241E-09-8.69954114E-14    2
-4.98606882E+03-7.00604665E+01-2.12213030E-01+6.87756030E-02-4.21067325E-05    3
+1.30061090E-08-1.60770046E-12+1.89801840E+03+3.18494469E+01+0.00000000E+00    4
C6H13-2                 C   6H  13    0    0G   300.000  5000.000 1396.000    51
+1.80640936E+01+2.85111833E-02-9.67861302E-06+1.49502045E-09-8.64303710E-14    2
-6.45433301E+03-6.70878929E+01+6.20068248E-01+6.16195063E-02-2.96980348E-05    3
+4.69998266E-09+3.13755723E-13+3.23741699E+02+2.92321681E+01+0.00000000E+00    4
C6H13-3                 C   6H  13    0    0G   300.000  5000.000 1396.000    51
+1.80640936E+01+2.85111833E-02-9.67861302E-06+1.49502045E-09-8.64303710E-14    2
-6.45433301E+03-6.70878929E+01+6.20068248E-01+6.16195063E-02-2.96980348E-05    3
+4.69998266E-09+3.13755723E-13+3.23741699E+02+2.92321681E+01+0.00000000E+00    4
C6H13OOH-1              C   6H  14O   2    0G   300.000  5000.000 1393.000    71
+2.45163599E+01+3.04358125E-02-1.04768961E-05+1.63358168E-09-9.50618695E-14    2
-4.15677013E+04-9.85011918E+01+3.76304221E-01+8.42019657E-02-5.55911124E-05    3
+1.86319290E-08-2.52819359E-12-3.29059850E+04+3.21031523E+01+0.00000000E+00    4
C6H13OOH-2              C   6H  14O   2    0G   300.000  5000.000 1401.000    71
+2.48832119E+01+2.96512073E-02-1.01015279E-05+1.56407586E-09-9.05729002E-14    2
-4.34204125E+04-1.01048943E+02+7.33867061E-01+8.64149041E-02-6.11174825E-05    3
+2.24268392E-08-3.36429856E-12-3.50923807E+04+2.84824773E+01+0.00000000E+00    4
C6H13OOH-3              C   6H  14O   2    0G   300.000  5000.000 1401.000    71
+2.48832119E+01+2.96512073E-02-1.01015279E-05+1.56407586E-09-9.05729002E-14    2
-4.34204125E+04-1.01048943E+02+7.33867061E-01+8.64149041E-02-6.11174825E-05    3
+2.24268392E-08-3.36429856E-12-3.50923807E+04+2.84824773E+01+0.00000000E+00    4
C6H13O2-1               C   6H  13O   2    0G   300.000  5000.000 1392.000    61
+2.31785440E+01+2.94255210E-02-1.01218190E-05+1.57735564E-09-9.17519123E-14    2
-2.41616714E+04-9.09398761E+01+1.05761492E+00+7.89345805E-02-5.23116185E-05    3
+1.79548180E-08-2.54740591E-12-1.62091180E+04+2.87209949E+01+0.00000000E+00    4
C6H13O2-2               C   6H  13O   2    0G   300.000  5000.000 1399.000    61
+2.34641557E+01+2.87030846E-02-9.76607754E-06+1.51070014E-09-8.74195382E-14    2
-2.59745219E+04-9.30010056E+01+1.59315499E+00+8.03858598E-02-5.68690473E-05    3
+2.12270568E-08-3.27992517E-12-1.84223008E+04+2.42747128E+01+0.00000000E+00    4
C6H13O2-3               C   6H  13O   2    0G   300.000  5000.000 1399.000    61
+2.34641557E+01+2.87030846E-02-9.76607754E-06+1.51070014E-09-8.74195382E-14    2
-2.59745219E+04-9.30010056E+01+1.59315499E+00+8.03858598E-02-5.68690473E-05    3
+2.12270568E-08-3.27992517E-12-1.84223008E+04+2.42747128E+01+0.00000000E+00    4
C6H13O-1                C   6H  13O   1    0G   300.000  5000.000 1396.000    51
+2.20928922E+01+2.79119481E-02-9.53349733E-06+1.47885354E-09-8.57536878E-14    2
-2.26216369E+04-8.78582845E+01+1.37476919E+00+7.09707741E-02-4.11061030E-05    3
+1.06839948E-08-8.50881624E-13-1.49531106E+04+2.52025044E+01+0.00000000E+00    4
C6H13O-2                C   6H  13O   1    0G   300.000  5000.000 1405.000    51
+2.18292052E+01+2.77008387E-02-9.36457645E-06+1.44248495E-09-8.32314882E-14    2
-2.43135941E+04-8.67680797E+01+1.53124348E+00+7.23874176E-02-4.54632890E-05    3
+1.39938106E-08-1.63272186E-12-1.70585882E+04+2.30983559E+01+0.00000000E+00    4
C6H13O-3                C   6H  13O   1    0G   300.000  5000.000 1405.000    51
+2.18292052E+01+2.77008387E-02-9.36457645E-06+1.44248495E-09-8.32314882E-14    2
-2.43135941E+04-8.67680797E+01+1.53124348E+00+7.23874176E-02-4.54632890E-05    3
+1.39938106E-08-1.63272186E-12-1.70585882E+04+2.30983559E+01+0.00000000E+00    4
C6H12OOH1-2             C   6H  13O   2    0G   300.000  5000.000 1392.000    71
+2.33958970E+01+2.87500915E-02-9.87479228E-06+1.53738184E-09-8.93686071E-14    2
-1.75002122E+04-8.93745541E+01+2.35234877E+00+7.42464378E-02-4.64307066E-05    3
+1.44953455E-08-1.79518968E-12-9.79913038E+03+2.49856776E+01+0.00000000E+00    4
C6H12OOH1-3             C   6H  13O   2    0G   300.000  5000.000 1396.000    71
+2.27895146E+01+2.89701974E-02-9.88728294E-06+1.53286753E-09-8.88486536E-14    2
-1.75428625E+04-8.54563755E+01+1.92496561E+00+7.24529009E-02-4.20779710E-05    3
+1.11647255E-08-9.59696372E-13-9.81550072E+03+2.83886795E+01+0.00000000E+00    4
C6H12OOH1-4             C   6H  13O   2    0G   300.000  5000.000 1396.000    71
+2.27895146E+01+2.89701974E-02-9.88728294E-06+1.53286753E-09-8.88486536E-14    2
-1.75428625E+04-8.54563755E+01+1.92496561E+00+7.24529009E-02-4.20779710E-05    3
+1.11647255E-08-9.59696372E-13-9.81550072E+03+2.83886795E+01+0.00000000E+00    4
C6H12OOH1-5             C   6H  13O   2    0G   300.000  5000.000 1396.000    71
+2.27895146E+01+2.89701974E-02-9.88728294E-06+1.53286753E-09-8.88486536E-14    2
-1.75428625E+04-8.54563755E+01+1.92496561E+00+7.24529009E-02-4.20779710E-05    3
+1.11647255E-08-9.59696372E-13-9.81550072E+03+2.83886795E+01+0.00000000E+00    4
C6H12OOH2-1             C   6H  13O   2    0G   300.000  5000.000 1401.000    71
+2.45762848E+01+2.74155943E-02-9.34192750E-06+1.44672243E-09-8.37892149E-14    2
-1.83935404E+04-9.65123105E+01+1.63351733E+00+8.14796740E-02-5.79995011E-05    3
+2.13418964E-08-3.19994195E-12-1.05064447E+04+2.64803283E+01+0.00000000E+00    4
C6H12OOH2-3             C   6H  13O   2    0G   300.000  5000.000 1400.000    71
+2.36864065E+01+2.80115990E-02-9.51112192E-06+1.46925773E-09-8.49419123E-14    2
-1.93109406E+04-9.14557581E+01+2.72663117E+00+7.64651999E-02-5.21833045E-05    3
+1.85187539E-08-2.69369864E-12-1.19891933E+04+2.12761646E+01+0.00000000E+00    4
C6H12OOH2-4             C   6H  13O   2    0G   300.000  5000.000 1408.000    71
+2.31606108E+01+2.80956105E-02-9.46369942E-06+1.45419355E-09-8.37638675E-14    2
-1.93834354E+04-8.79850394E+01+2.26007590E+00+7.48358213E-02-4.80375241E-05    3
+1.52775741E-08-1.87091068E-12-1.19995231E+04+2.48618430E+01+0.00000000E+00    4
C6H12OOH2-5             C   6H  13O   2    0G   300.000  5000.000 1408.000    71
+2.31606108E+01+2.80956105E-02-9.46369942E-06+1.45419355E-09-8.37638675E-14    2
-1.93834354E+04-8.79850394E+01+2.26007590E+00+7.48358213E-02-4.80375241E-05    3
+1.52775741E-08-1.87091068E-12-1.19995231E+04+2.48618430E+01+0.00000000E+00    4
C6H12OOH2-6             C   6H  13O   2    0G   300.000  5000.000 1402.000    71
+2.43039070E+01+2.76074809E-02-9.39913372E-06+1.45469578E-09-8.42141472E-14    2
-1.82854496E+04-9.51106853E+01+1.09455724E+00+8.29967617E-02-6.01254476E-05    3
+2.26497954E-08-3.48706819E-12-1.03716865E+04+2.90715700E+01+0.00000000E+00    4
C6H12OOH3-1             C   6H  13O   2    0G   300.000  5000.000 1402.000    71
+2.43039070E+01+2.76074809E-02-9.39913372E-06+1.45469578E-09-8.42141472E-14    2
-1.82854496E+04-9.51106853E+01+1.09455724E+00+8.29967617E-02-6.01254476E-05    3
+2.26497954E-08-3.48706819E-12-1.03716865E+04+2.90715700E+01+0.00000000E+00    4
C6H12OOH3-2             C   6H  13O   2    0G   300.000  5000.000 1400.000    71
+2.36864065E+01+2.80115990E-02-9.51112192E-06+1.46925773E-09-8.49419123E-14    2
-1.93109406E+04-9.14557581E+01+2.72663117E+00+7.64651999E-02-5.21833045E-05    3
+1.85187539E-08-2.69369864E-12-1.19891933E+04+2.12761646E+01+0.00000000E+00    4
C6H12OOH3-4             C   6H  13O   2    0G   300.000  5000.000 1400.000    71
+2.36864065E+01+2.80115990E-02-9.51112192E-06+1.46925773E-09-8.49419123E-14    2
-1.93109406E+04-9.14557581E+01+2.72663117E+00+7.64651999E-02-5.21833045E-05    3
+1.85187539E-08-2.69369864E-12-1.19891933E+04+2.12761646E+01+0.00000000E+00    4
C6H12OOH3-5             C   6H  13O   2    0G   300.000  5000.000 1408.000    71
+2.31606108E+01+2.80956105E-02-9.46369942E-06+1.45419355E-09-8.37638675E-14    2
-1.93834354E+04-8.79850394E+01+2.26007590E+00+7.48358213E-02-4.80375241E-05    3
+1.52775741E-08-1.87091068E-12-1.19995231E+04+2.48618430E+01+0.00000000E+00    4
C6H12OOH3-6             C   6H  13O   2    0G   300.000  5000.000 1402.000    71
+2.43039070E+01+2.76074809E-02-9.39913372E-06+1.45469578E-09-8.42141472E-14    2
-1.82854496E+04-9.51106853E+01+1.09455724E+00+8.29967617E-02-6.01254476E-05    3
+2.26497954E-08-3.48706819E-12-1.03716865E+04+2.90715700E+01+0.00000000E+00    4
C6H12O1-2               C   6H  12O   1    0G   300.000  5000.000 1418.000    41
+2.09805167E+01+2.61456832E-02-8.79805046E-06+1.35121022E-09-7.78107305E-14    2
-2.91366825E+04-8.58639749E+01-5.27479473E+00+9.15832630E-02-7.09194990E-05    3
+2.79461610E-08-4.39482049E-12-2.05857903E+04+5.34224762E+01+0.00000000E+00    4
C6H12O1-3               C   6H  12O   1    0G   300.000  5000.000 1412.000    31
+1.99712630E+01+2.75739130E-02-9.32003684E-06+1.43550676E-09-8.28258579E-14    2
-2.99062932E+04-8.20867887E+01-8.93042069E+00+1.02982605E-01-8.53638224E-05    3
+3.63896486E-08-6.21235185E-12-2.07664357E+04+7.01497676E+01+0.00000000E+00    4
C6H12O1-4               C   6H  12O   1    0G   300.000  5000.000 1451.000    21
+1.87967925E+01+2.75535527E-02-9.00773471E-06+1.35601108E-09-7.69845934E-14    2
-3.93246166E+04-7.58383918E+01-8.12435380E+00+9.70640114E-02-7.69405734E-05    3
+3.10474493E-08-4.95396033E-12-3.08886808E+04+6.59704356E+01+0.00000000E+00    4
C6H12O1-5               C   6H  12O   1    0G   300.000  5000.000 1411.000    11
+1.99284959E+01+2.86967410E-02-9.76084126E-06+1.50996782E-09-8.73930262E-14    2
-4.25348728E+04-8.86574195E+01-1.13294962E+01+1.08590522E-01-8.83887484E-05    3
+3.67290337E-08-6.10865223E-12-3.24988594E+04+7.65557826E+01+0.00000000E+00    4
C6H12O2-3               C   6H  12O   1    0G   300.000  5000.000 1425.000    41
+2.14267419E+01+2.53570884E-02-8.43894210E-06+1.28635266E-09-7.36861092E-14    2
-3.11276934E+04-8.88992853E+01-5.25994961E+00+9.41384839E-02-7.60798059E-05    3
+3.12814710E-08-5.11045005E-12-2.26926336E+04+5.18211467E+01+0.00000000E+00    4
C6H12O2-4               C   6H  12O   1    0G   300.000  5000.000 1417.000    31
+2.02636052E+01+2.68979324E-02-8.99457950E-06+1.37527090E-09-7.89420963E-14    2
-3.18212913E+04-8.42025816E+01-8.71729383E+00+1.04644598E-01-8.94323784E-05    3
+3.91535754E-08-6.81619305E-12-2.29012647E+04+6.76413269E+01+0.00000000E+00    4
C6H12O2-5               C   6H  12O   1    0G   300.000  5000.000 1418.000    21
+1.96691261E+01+2.77995312E-02-9.30042882E-06+1.42255648E-09-8.16795227E-14    2
-4.19335698E+04-8.31528662E+01-1.07496328E+01+1.08968762E-01-9.26948775E-05    3
+4.02824223E-08-6.95618656E-12-3.25413826E+04+7.63557140E+01+0.00000000E+00    4
C6H12O3-4               C   6H  12O   1    0G   300.000  5000.000 1425.000    41
+2.14267419E+01+2.53570884E-02-8.43894210E-06+1.28635266E-09-7.36861092E-14    2
-3.11276934E+04-8.95887669E+01-5.25994961E+00+9.41384839E-02-7.60798059E-05    3
+3.12814710E-08-5.11045005E-12-2.26926336E+04+5.11316651E+01+0.00000000E+00    4
C6H12OOH1-2O2           C   6H  13O   4    0G   300.000  5000.000 1394.000    81
+3.04683025E+01+2.77522708E-02-9.61137583E-06+1.50516303E-09-8.78680262E-14    2
-3.83461529E+04-1.25345284E+02+2.62680845E+00+8.94856642E-02-5.98279275E-05    3
+1.91011928E-08-2.28528990E-12-2.84709479E+04+2.51462108E+01+0.00000000E+00    4
C6H12OOH1-3O2           C   6H  13O   4    0G   300.000  5000.000 1394.000    81
+3.04683025E+01+2.77522708E-02-9.61137583E-06+1.50516303E-09-8.78680262E-14    2
-3.83461529E+04-1.25345284E+02+2.62680845E+00+8.94856642E-02-5.98279275E-05    3
+1.91011928E-08-2.28528990E-12-2.84709479E+04+2.51462108E+01+0.00000000E+00    4
C6H12OOH1-4O2           C   6H  13O   4    0G   300.000  5000.000 1394.000    81
+3.04683025E+01+2.77522708E-02-9.61137583E-06+1.50516303E-09-8.78680262E-14    2
-3.83461529E+04-1.25345284E+02+2.62680845E+00+8.94856642E-02-5.98279275E-05    3
+1.91011928E-08-2.28528990E-12-2.84709479E+04+2.51462108E+01+0.00000000E+00    4
C6H12OOH1-5O2           C   6H  13O   4    0G   300.000  5000.000 1394.000    81
+3.04683025E+01+2.77522708E-02-9.61137583E-06+1.50516303E-09-8.78680262E-14    2
-3.83461529E+04-1.25345284E+02+2.62680845E+00+8.94856642E-02-5.98279275E-05    3
+1.91011928E-08-2.28528990E-12-2.84709479E+04+2.51462108E+01+0.00000000E+00    4
C6H12OOH2-1O2           C   6H  13O   4    0G   300.000  5000.000 1394.000    81
+3.04683025E+01+2.77522708E-02-9.61137583E-06+1.50516303E-09-8.78680262E-14    2
-3.83461529E+04-1.25345284E+02+2.62680845E+00+8.94856642E-02-5.98279275E-05    3
+1.91011928E-08-2.28528990E-12-2.84709479E+04+2.51462108E+01+0.00000000E+00    4
C6H12OOH2-3O2           C   6H  13O   4    0G   300.000  5000.000 1403.000    81
+2.83590321E+01+2.87735842E-02-9.78879765E-06+1.51428335E-09-8.76360651E-14    2
-3.91336282E+04-1.13425601E+02+2.53306668E+00+9.21554288E-02-6.98231363E-05    3
+2.75462625E-08-4.42827896E-12-3.05121822E+04+2.41208096E+01+0.00000000E+00    4
C6H12OOH2-4O2           C   6H  13O   4    0G   300.000  5000.000 1403.000    81
+2.83590321E+01+2.87735842E-02-9.78879765E-06+1.51428335E-09-8.76360651E-14    2
-3.91336282E+04-1.13425601E+02+2.53306668E+00+9.21554288E-02-6.98231363E-05    3
+2.75462625E-08-4.42827896E-12-3.05121822E+04+2.41208096E+01+0.00000000E+00    4
C6H12OOH2-5O2           C   6H  13O   4    0G   300.000  5000.000 1403.000    81
+2.83590321E+01+2.87735842E-02-9.78879765E-06+1.51428335E-09-8.76360651E-14    2
-3.91336282E+04-1.13425601E+02+2.53306668E+00+9.21554288E-02-6.98231363E-05    3
+2.75462625E-08-4.42827896E-12-3.05121822E+04+2.41208096E+01+0.00000000E+00    4
C6H12OOH2-6O2           C   6H  13O   4    0G   300.000  5000.000 1394.000    81
+3.04683025E+01+2.77522708E-02-9.61137583E-06+1.50516303E-09-8.78680262E-14    2
-3.83461529E+04-1.25345284E+02+2.62680845E+00+8.94856642E-02-5.98279275E-05    3
+1.91011928E-08-2.28528990E-12-2.84709479E+04+2.51462108E+01+0.00000000E+00    4
C6H12OOH3-1O2           C   6H  13O   4    0G   300.000  5000.000 1394.000    81
+3.04683025E+01+2.77522708E-02-9.61137583E-06+1.50516303E-09-8.78680262E-14    2
-3.83461529E+04-1.25345284E+02+2.62680845E+00+8.94856642E-02-5.98279275E-05    3
+1.91011928E-08-2.28528990E-12-2.84709479E+04+2.51462108E+01+0.00000000E+00    4
C6H12OOH3-2O2           C   6H  13O   4    0G   300.000  5000.000 1403.000    81
+2.83590321E+01+2.87735842E-02-9.78879765E-06+1.51428335E-09-8.76360651E-14    2
-3.91336282E+04-1.13425601E+02+2.53306668E+00+9.21554288E-02-6.98231363E-05    3
+2.75462625E-08-4.42827896E-12-3.05121822E+04+2.41208096E+01+0.00000000E+00    4
C6H12OOH3-4O2           C   6H  13O   4    0G   300.000  5000.000 1403.000    81
+2.83590321E+01+2.87735842E-02-9.78879765E-06+1.51428335E-09-8.76360651E-14    2
-3.91336282E+04-1.13425601E+02+2.53306668E+00+9.21554288E-02-6.98231363E-05    3
+2.75462625E-08-4.42827896E-12-3.05121822E+04+2.41208096E+01+0.00000000E+00    4
C6H12OOH3-5O2           C   6H  13O   4    0G   300.000  5000.000 1403.000    81
+2.83590321E+01+2.87735842E-02-9.78879765E-06+1.51428335E-09-8.76360651E-14    2
-3.91336282E+04-1.13425601E+02+2.53306668E+00+9.21554288E-02-6.98231363E-05    3
+2.75462625E-08-4.42827896E-12-3.05121822E+04+2.41208096E+01+0.00000000E+00    4
C6H12OOH3-6O2           C   6H  13O   4    0G   300.000  5000.000 1394.000    81
+3.04683025E+01+2.77522708E-02-9.61137583E-06+1.50516303E-09-8.78680262E-14    2
-3.83461529E+04-1.25345284E+02+2.62680845E+00+8.94856642E-02-5.98279275E-05    3
+1.91011928E-08-2.28528990E-12-2.84709479E+04+2.51462108E+01+0.00000000E+00    4
C6H11-1D3OOH            C   6H  12O   2    0G   300.000  5000.000 1393.000    61
+2.59035094E+01+2.42696112E-02-8.29035467E-06+1.28689728E-09-7.46830616E-14    2
-2.68476823E+04-1.07452182E+02-2.31977696E+00+9.52241599E-02-7.73053497E-05    3
+3.20512066E-08-5.34750057E-12-1.76191545E+04+4.22269905E+01+0.00000000E+00    4
C6H11-1D4OOH            C   6H  12O   2    0G   300.000  5000.000 1401.000    61
+2.29270511E+01+2.66225664E-02-9.05133554E-06+1.39947254E-09-8.09578355E-14    2
-2.71948840E+04-8.94129595E+01+1.13416759E+00+7.94193160E-02-5.85260848E-05    3
+2.26979408E-08-3.62009744E-12-1.98209376E+04+2.69474429E+01+0.00000000E+00    4
C6H11-1D5OOH            C   6H  12O   2    0G   300.000  5000.000 1401.000    61
+2.29270511E+01+2.66225664E-02-9.05133554E-06+1.39947254E-09-8.09578355E-14    2
-2.71948840E+04-8.94129595E+01+1.13416759E+00+7.94193160E-02-5.85260848E-05    3
+2.26979408E-08-3.62009744E-12-1.98209376E+04+2.69474429E+01+0.00000000E+00    4
C6H11-1D6OOH            C   6H  12O   2    0G   300.000  5000.000 1393.000    61
+2.26383519E+01+2.73757543E-02-9.42397309E-06+1.46942591E-09-8.55091451E-14    2
-2.53967947E+04-8.73725472E+01+6.48701799E-01+7.76335542E-02-5.34143826E-05    3
+1.90936716E-08-2.82021629E-12-1.76120903E+04+3.11812799E+01+0.00000000E+00    4
C6H11-2D1OOH            C   6H  12O   2    0G   300.000  5000.000 1385.000    61
+2.43428219E+01+2.60142938E-02-8.97949936E-06+1.40314527E-09-8.17901261E-14    2
-2.57267860E+04-9.65749831E+01+2.11692928E-01+8.23288253E-02-5.97664416E-05    3
+2.25592257E-08-3.51959321E-12-1.72986603E+04+3.31182384E+01+0.00000000E+00    4
C6H11-2D4OOH            C   6H  12O   2    0G   300.000  5000.000 1392.000    61
+2.53272397E+01+2.47729296E-02-8.46596932E-06+1.31443483E-09-7.62890280E-14    2
-2.79852809E+04-1.04859678E+02-1.46245581E+00+9.02938420E-02-7.01570906E-05    3
+2.78745585E-08-4.47562215E-12-1.90395758E+04+3.78704689E+01+0.00000000E+00    4
C6H11-2D5OOH            C   6H  12O   2    0G   300.000  5000.000 1399.000    61
+2.25048513E+01+2.69114345E-02-9.13654120E-06+1.41134534E-09-8.15937722E-14    2
-2.83951897E+04-8.76985785E+01+1.81623661E+00+7.52045876E-02-5.22511183E-05    3
+1.89442291E-08-2.82183511E-12-2.12139988E+04+2.34113083E+01+0.00000000E+00    4
C6H11-2D6OOH            C   6H  12O   2    0G   300.000  5000.000 1390.000    61
+2.21518946E+01+2.77388788E-02-9.53838077E-06+1.48617108E-09-8.64396575E-14    2
-2.65647544E+04-8.52712241E+01+1.51940041E+00+7.26401571E-02-4.60784955E-05    3
+1.47295637E-08-1.89409854E-12-1.90350093E+04+2.67655882E+01+0.00000000E+00    4
C6H11-3D1OOH            C   6H  12O   2    0G   300.000  5000.000 1390.000    61
+2.18169743E+01+2.80152259E-02-9.63205183E-06+1.50063123E-09-8.72754508E-14    2
-2.64614918E+04-8.35297001E+01+1.17006930E+00+7.27400593E-02-4.57945723E-05    3
+1.44941072E-08-1.84089055E-12-1.89021358E+04+2.86651787E+01+0.00000000E+00    4
C6H11-3D2OOH            C   6H  12O   2    0G   300.000  5000.000 1391.000    61
+2.50642842E+01+2.49351789E-02-8.51039657E-06+1.32031801E-09-7.65936140E-14    2
-2.79114429E+04-1.03524314E+02-1.79725520E+00+9.02776158E-02-6.96160763E-05    3
+2.74275414E-08-4.36716320E-12-1.89077528E+04+3.97122202E+01+0.00000000E+00    4
C6H11Q12-3              C   6H  13O   4    0G   300.000  5000.000 1394.000    91
+2.78943291E+01+2.92847808E-02-1.00847792E-05+1.57294057E-09-9.15554523E-14    2
-3.05839622E+04-1.07701979E+02+2.99684347E+00+8.60938560E-02-5.92978062E-05    3
+2.08719630E-08-2.98876240E-12-2.18052539E+04+2.64874463E+01+0.00000000E+00    4
C6H11Q12-4              C   6H  13O   4    0G   300.000  5000.000 1409.000    91
+2.80581380E+01+2.85464861E-02-9.69832158E-06+1.49895066E-09-8.66960196E-14    2
-3.05545861E+04-1.07396273E+02+3.80954684E+00+8.47207481E-02-5.85351924E-05    3
+2.03764845E-08-2.81456479E-12-2.21836150E+04+2.28354127E+01+0.00000000E+00    4
C6H11Q12-5              C   6H  13O   4    0G   300.000  5000.000 1409.000    91
+2.80581380E+01+2.85464861E-02-9.69832158E-06+1.49895066E-09-8.66960196E-14    2
-3.05545861E+04-1.07396273E+02+3.80954684E+00+8.47207481E-02-5.85351924E-05    3
+2.03764845E-08-2.81456479E-12-2.21836150E+04+2.28354127E+01+0.00000000E+00    4
C6H11Q12-6              C   6H  13O   4    0G   300.000  5000.000 1396.000    91
+3.09468859E+01+2.69623754E-02-9.34843940E-06+1.46514666E-09-8.55805589E-14    2
-3.04867475E+04-1.25320374E+02+2.20320858E+00+9.20185664E-02-6.38825199E-05    3
+2.14499236E-08-2.76271950E-12-2.04338777E+04+2.95618135E+01+0.00000000E+00    4
C6H11Q13-2              C   6H  13O   4    0G   300.000  5000.000 1394.000    91
+2.78943291E+01+2.92847808E-02-1.00847792E-05+1.57294057E-09-9.15554523E-14    2
-3.05839622E+04-1.07701979E+02+2.99684347E+00+8.60938560E-02-5.92978062E-05    3
+2.08719630E-08-2.98876240E-12-2.18052539E+04+2.64874463E+01+0.00000000E+00    4
C6H11Q13-4              C   6H  13O   4    0G   300.000  5000.000 1394.000    91
+2.78943291E+01+2.92847808E-02-1.00847792E-05+1.57294057E-09-9.15554523E-14    2
-3.05839622E+04-1.07701979E+02+2.99684347E+00+8.60938560E-02-5.92978062E-05    3
+2.08719630E-08-2.98876240E-12-2.18052539E+04+2.64874463E+01+0.00000000E+00    4
C6H11Q13-5              C   6H  13O   4    0G   300.000  5000.000 1409.000    91
+2.80581380E+01+2.85464861E-02-9.69832158E-06+1.49895066E-09-8.66960196E-14    2
-3.05545861E+04-1.07396273E+02+3.80954684E+00+8.47207481E-02-5.85351924E-05    3
+2.03764845E-08-2.81456479E-12-2.21836150E+04+2.28354127E+01+0.00000000E+00    4
C6H11Q13-6              C   6H  13O   4    0G   300.000  5000.000 1396.000    91
+3.09468859E+01+2.69623754E-02-9.34843940E-06+1.46514666E-09-8.55805589E-14    2
-3.04867475E+04-1.25320374E+02+2.20320858E+00+9.20185664E-02-6.38825199E-05    3
+2.14499236E-08-2.76271950E-12-2.04338777E+04+2.95618135E+01+0.00000000E+00    4
C6H11Q14-2              C   6H  13O   4    0G   300.000  5000.000 1394.000    91
+2.78943291E+01+2.92847808E-02-1.00847792E-05+1.57294057E-09-9.15554523E-14    2
-3.05839622E+04-1.07701979E+02+2.99684347E+00+8.60938560E-02-5.92978062E-05    3
+2.08719630E-08-2.98876240E-12-2.18052539E+04+2.64874463E+01+0.00000000E+00    4
C6H11Q14-3              C   6H  13O   4    0G   300.000  5000.000 1394.000    91
+2.78943291E+01+2.92847808E-02-1.00847792E-05+1.57294057E-09-9.15554523E-14    2
-3.05839622E+04-1.07701979E+02+2.99684347E+00+8.60938560E-02-5.92978062E-05    3
+2.08719630E-08-2.98876240E-12-2.18052539E+04+2.64874463E+01+0.00000000E+00    4
C6H11Q14-5              C   6H  13O   4    0G   300.000  5000.000 1394.000    91
+2.78943291E+01+2.92847808E-02-1.00847792E-05+1.57294057E-09-9.15554523E-14    2
-3.05839622E+04-1.07701979E+02+2.99684347E+00+8.60938560E-02-5.92978062E-05    3
+2.08719630E-08-2.98876240E-12-2.18052539E+04+2.64874463E+01+0.00000000E+00    4
C6H11Q14-6              C   6H  13O   4    0G   300.000  5000.000 1396.000    91
+3.09468859E+01+2.69623754E-02-9.34843940E-06+1.46514666E-09-8.55805589E-14    2
-3.04867475E+04-1.25320374E+02+2.20320858E+00+9.20185664E-02-6.38825199E-05    3
+2.14499236E-08-2.76271950E-12-2.04338777E+04+2.95618135E+01+0.00000000E+00    4
C6H11Q15-2              C   6H  13O   4    0G   300.000  5000.000 1394.000    91
+2.78943291E+01+2.92847808E-02-1.00847792E-05+1.57294057E-09-9.15554523E-14    2
-3.05839622E+04-1.07701979E+02+2.99684347E+00+8.60938560E-02-5.92978062E-05    3
+2.08719630E-08-2.98876240E-12-2.18052539E+04+2.64874463E+01+0.00000000E+00    4
C6H11Q15-3              C   6H  13O   4    0G   300.000  5000.000 1409.000    91
+2.80581380E+01+2.85464861E-02-9.69832158E-06+1.49895066E-09-8.66960196E-14    2
-3.05545861E+04-1.07396273E+02+3.80954684E+00+8.47207481E-02-5.85351924E-05    3
+2.03764845E-08-2.81456479E-12-2.21836150E+04+2.28354127E+01+0.00000000E+00    4
C6H11Q15-4              C   6H  13O   4    0G   300.000  5000.000 1394.000    91
+2.78943291E+01+2.92847808E-02-1.00847792E-05+1.57294057E-09-9.15554523E-14    2
-3.05839622E+04-1.07701979E+02+2.99684347E+00+8.60938560E-02-5.92978062E-05    3
+2.08719630E-08-2.98876240E-12-2.18052539E+04+2.64874463E+01+0.00000000E+00    4
C6H11Q15-6              C   6H  13O   4    0G   300.000  5000.000 1396.000    91
+2.82883945E+01+2.89369583E-02-9.96190727E-06+1.55346138E-09-9.04091590E-14    2
-2.93711746E+04-1.09680591E+02+2.12435546E+00+9.08091150E-02-6.62026612E-05    3
+2.49559670E-08-3.84884889E-12-2.03676921E+04+3.05566985E+01+0.00000000E+00    4
C6H11Q23-1              C   6H  13O   4    0G   300.000  5000.000 1402.000    91
+2.87206101E+01+2.81926003E-02-9.62199118E-06+1.49176614E-09-8.64680578E-14    2
-3.13085620E+04-1.12729880E+02+2.50274303E+00+9.23699697E-02-7.01978035E-05    3
+2.76525328E-08-4.43054874E-12-2.25427916E+04+2.69579667E+01+0.00000000E+00    4
C6H11Q23-4              C   6H  13O   4    0G   300.000  5000.000 1400.000    91
+2.83307086E+01+2.85436428E-02-9.74746596E-06+1.51180692E-09-8.76533346E-14    2
-3.25271405E+04-1.10789659E+02+3.37103808E+00+8.76299651E-02-6.32127378E-05    3
+2.35062741E-08-3.55550322E-12-2.39785960E+04+2.29119049E+01+0.00000000E+00    4
C6H11Q23-5              C   6H  13O   4    0G   300.000  5000.000 1421.000    91
+2.84438571E+01+2.76525438E-02-9.26702496E-06+1.41900244E-09-8.15353368E-14    2
-3.24103661E+04-1.10029025E+02+4.01277430E+00+8.75230514E-02-6.49830548E-05    3
+2.47375697E-08-3.77261053E-12-2.43431110E+04+1.99545556E+01+0.00000000E+00    4
C6H11Q23-6              C   6H  13O   4    0G   300.000  5000.000 1403.000    91
+2.86807869E+01+2.81353066E-02-9.58211151E-06+1.48344887E-09-8.58991774E-14    2
-3.12397030E+04-1.12551544E+02+2.07300290E+00+9.43156884E-02-7.32191610E-05    3
+2.95085081E-08-4.82851589E-12-2.24527685E+04+2.88342959E+01+0.00000000E+00    4
C6H11Q24-1              C   6H  13O   4    0G   300.000  5000.000 1402.000    91
+2.87206101E+01+2.81926003E-02-9.62199118E-06+1.49176614E-09-8.64680578E-14    2
-3.13085620E+04-1.12729880E+02+2.50274303E+00+9.23699697E-02-7.01978035E-05    3
+2.76525328E-08-4.43054874E-12-2.25427916E+04+2.69579667E+01+0.00000000E+00    4
C6H11Q24-3              C   6H  13O   4    0G   300.000  5000.000 1400.000    91
+2.83307086E+01+2.85436428E-02-9.74746596E-06+1.51180692E-09-8.76533346E-14    2
-3.25271405E+04-1.10789659E+02+3.37103808E+00+8.76299651E-02-6.32127378E-05    3
+2.35062741E-08-3.55550322E-12-2.39785960E+04+2.29119049E+01+0.00000000E+00    4
C6H11Q24-5              C   6H  13O   4    0G   300.000  5000.000 1400.000    91
+2.83307086E+01+2.85436428E-02-9.74746596E-06+1.51180692E-09-8.76533346E-14    2
-3.25271405E+04-1.10789659E+02+3.37103808E+00+8.76299651E-02-6.32127378E-05    3
+2.35062741E-08-3.55550322E-12-2.39785960E+04+2.29119049E+01+0.00000000E+00    4
C6H11Q24-6              C   6H  13O   4    0G   300.000  5000.000 1403.000    91
+2.86807869E+01+2.81353066E-02-9.58211151E-06+1.48344887E-09-8.58991774E-14    2
-3.12397030E+04-1.12551544E+02+2.07300290E+00+9.43156884E-02-7.32191610E-05    3
+2.95085081E-08-4.82851589E-12-2.24527685E+04+2.88342959E+01+0.00000000E+00    4
C6H11Q25-1              C   6H  13O   4    0G   300.000  5000.000 1402.000    91
+2.87206101E+01+2.81926003E-02-9.62199118E-06+1.49176614E-09-8.64680578E-14    2
-3.13085620E+04-1.12729880E+02+2.50274303E+00+9.23699697E-02-7.01978035E-05    3
+2.76525328E-08-4.43054874E-12-2.25427916E+04+2.69579667E+01+0.00000000E+00    4
C6H11Q25-3              C   6H  13O   4    0G   300.000  5000.000 1400.000    91
+2.83307086E+01+2.85436428E-02-9.74746596E-06+1.51180692E-09-8.76533346E-14    2
-3.25271405E+04-1.10789659E+02+3.37103808E+00+8.76299651E-02-6.32127378E-05    3
+2.35062741E-08-3.55550322E-12-2.39785960E+04+2.29119049E+01+0.00000000E+00    4
C6H11Q34-1              C   6H  13O   4    0G   300.000  5000.000 1403.000    91
+2.86807869E+01+2.81353066E-02-9.58211151E-06+1.48344887E-09-8.58991774E-14    2
-3.12397030E+04-1.12551544E+02+2.07300290E+00+9.43156884E-02-7.32191610E-05    3
+2.95085081E-08-4.82851589E-12-2.24527685E+04+2.88342959E+01+0.00000000E+00    4
C6H11Q34-2              C   6H  13O   4    0G   300.000  5000.000 1400.000    91
+2.83307086E+01+2.85436428E-02-9.74746596E-06+1.51180692E-09-8.76533346E-14    2
-3.25271405E+04-1.10789659E+02+3.37103808E+00+8.76299651E-02-6.32127378E-05    3
+2.35062741E-08-3.55550322E-12-2.39785960E+04+2.29119049E+01+0.00000000E+00    4
C6KET12                 C   6H  12O   3    0G   300.000  5000.000 1387.000    71
+2.90256185E+01+2.40820489E-02-8.30639705E-06+1.29822444E-09-7.57124082E-14    2
-5.32782165E+04-1.19864821E+02-1.70742664E+00+9.97939251E-02-8.01901862E-05    3
+3.25346440E-08-5.30122784E-12-4.30784665E+04+4.36695548E+01+0.00000000E+00    4
C6KET13                 C   6H  12O   3    0G   300.000  5000.000 1403.000    71
+2.58825405E+01+2.62029247E-02-8.90539787E-06+1.37704650E-09-7.96812443E-14    2
-5.34388150E+04-1.02769588E+02+2.70686236E+00+7.86587312E-02-5.28474860E-05    3
+1.74402371E-08-2.21798402E-12-4.53342182E+04+2.21065759E+01+0.00000000E+00    4
C6KET14                 C   6H  12O   3    0G   300.000  5000.000 1403.000    71
+2.58825405E+01+2.62029247E-02-8.90539787E-06+1.37704650E-09-7.96812443E-14    2
-5.34388150E+04-1.02769588E+02+2.70686236E+00+7.86587312E-02-5.28474860E-05    3
+1.74402371E-08-2.21798402E-12-4.53342182E+04+2.21065759E+01+0.00000000E+00    4
C6KET15                 C   6H  12O   3    0G   300.000  5000.000 1403.000    71
+2.58825405E+01+2.62029247E-02-8.90539787E-06+1.37704650E-09-7.96812443E-14    2
-5.34388150E+04-1.02769588E+02+2.70686236E+00+7.86587312E-02-5.28474860E-05    3
+1.74402371E-08-2.21798402E-12-4.53342182E+04+2.21065759E+01+0.00000000E+00    4
C6KET21                 C   6H  12O   3    0G   300.000  5000.000 1389.000    71
+2.79607714E+01+2.42379297E-02-8.20343155E-06+1.26648645E-09-7.32501537E-14    2
-5.43857540E+04-1.13016914E+02-5.14482555E-01+9.21784846E-02-6.94513152E-05    3
+2.60396658E-08-3.86537916E-12-4.47938808E+04+3.91532333E+01+0.00000000E+00    4
C6KET23                 C   6H  12O   3    0G   300.000  5000.000 1389.000    71
+2.77518536E+01+2.44228814E-02-8.26691484E-06+1.27620900E-09-7.38039402E-14    2
-5.63515030E+04-1.12222879E+02-8.86325259E-01+9.56932379E-02-7.66622031E-05    3
+3.13003623E-08-5.14052764E-12-4.69292576E+04+3.98915047E+01+0.00000000E+00    4
C6KET24                 C   6H  12O   3    0G   300.000  5000.000 1410.000    71
+2.45827447E+01+2.65291227E-02-8.85055847E-06+1.35140650E-09-7.75076694E-14    2
-5.64887218E+04-9.49507504E+01+3.38656723E+00+7.51931934E-02-5.03122375E-05    3
+1.68156568E-08-2.18752991E-12-4.91634551E+04+1.89837711E+01+0.00000000E+00    4
C6KET25                 C   6H  12O   3    0G   300.000  5000.000 1410.000    71
+2.45827447E+01+2.65291227E-02-8.85055847E-06+1.35140650E-09-7.75076694E-14    2
-5.64887218E+04-9.49507504E+01+3.38656723E+00+7.51931934E-02-5.03122375E-05    3
+1.68156568E-08-2.18752991E-12-4.91634551E+04+1.89837711E+01+0.00000000E+00    4
C6KET26                 C   6H  12O   3    0G   300.000  5000.000 1396.000    71
+2.41192811E+01+2.75685546E-02-9.34714604E-06+1.44293337E-09-8.33930684E-14    2
-5.46176520E+04-9.19195513E+01+2.91522244E+00+7.34293670E-02-4.53418223E-05    3
+1.33776385E-08-1.43669218E-12-4.69588500E+04+2.31405529E+01+0.00000000E+00    4
C6KET31                 C   6H  12O   3    0G   300.000  5000.000 1513.000    71
+2.47427707E+01+2.65724465E-02-8.91511787E-06+1.36741583E-09-7.87033305E-14    2
-5.49929590E+04-9.61506620E+01+3.68645338E+00+6.79151683E-02-3.49002426E-05    3
+5.86626515E-09+3.80680692E-13-4.70773283E+04+1.94153944E+01+0.00000000E+00    4
C6KET32                 C   6H  12O   3    0G   300.000  5000.000 1388.000    71
+2.78409221E+01+2.43352401E-02-8.23613901E-06+1.27151170E-09-7.35397855E-14    2
-5.65357668E+04-1.13496792E+02-3.40401334E-02+9.00007504E-02-6.64122175E-05    3
+2.42781825E-08-3.49817449E-12-4.70631692E+04+3.57622287E+01+0.00000000E+00    4
C6KET34                 C   6H  12O   3    0G   300.000  5000.000 1388.000    71
+2.78409221E+01+2.43352401E-02-8.23613901E-06+1.27151170E-09-7.35397855E-14    2
-5.65357668E+04-1.13496792E+02-3.40401334E-02+9.00007504E-02-6.64122175E-05    3
+2.42781825E-08-3.49817449E-12-4.70631692E+04+3.57622287E+01+0.00000000E+00    4
C6KET35                 C   6H  12O   3    0G   300.000  5000.000 1422.000    71
+2.52008823E+01+2.55867980E-02-8.44943107E-06+1.28209867E-09-7.32384055E-14    2
-5.68781816E+04-9.91884828E+01+4.11000703E+00+6.98568662E-02-4.01291482E-05    3
+9.49599829E-09-4.21088500E-13-4.92736613E+04+1.54877708E+01+0.00000000E+00    4
C6KET36                 C   6H  12O   3    0G   300.000  5000.000 1513.000    71
+2.47427707E+01+2.65724465E-02-8.91511787E-06+1.36741583E-09-7.87033305E-14    2
-5.49929590E+04-9.61506620E+01+3.68645338E+00+6.79151683E-02-3.49002426E-05    3
+5.86626515E-09+3.80680692E-13-4.70773283E+04+1.94153944E+01+0.00000000E+00    4
C6H11O12-3OOH           C   6H  12O   3    0G   300.000  5000.000 1432.000    61
+2.74037429E+01+2.47674765E-02-8.29487594E-06+1.27052501E-09-7.30489658E-14    2
-4.27151891E+04-1.14645759E+02-2.27599349E+00+9.86141518E-02-7.74723381E-05    3
+3.01376954E-08-4.58669108E-12-3.31277592E+04+4.27007503E+01+0.00000000E+00    4
C6H11O12-4OOH           C   6H  12O   3    0G   300.000  5000.000 1432.000    61
+2.74037429E+01+2.47674765E-02-8.29487594E-06+1.27052501E-09-7.30489658E-14    2
-4.27151891E+04-1.14645759E+02-2.27599349E+00+9.86141518E-02-7.74723381E-05    3
+3.01376954E-08-4.58669108E-12-3.31277592E+04+4.27007503E+01+0.00000000E+00    4
C6H11O12-5OOH           C   6H  12O   3    0G   300.000  5000.000 1432.000    61
+2.74037429E+01+2.47674765E-02-8.29487594E-06+1.27052501E-09-7.30489658E-14    2
-4.27151891E+04-1.14645759E+02-2.27599349E+00+9.86141518E-02-7.74723381E-05    3
+3.01376954E-08-4.58669108E-12-3.31277592E+04+4.27007503E+01+0.00000000E+00    4
C6H11O12-6OOH           C   6H  12O   3    0G   300.000  5000.000 1418.000    61
+2.64398182E+01+2.60261489E-02-8.81968488E-06+1.36137474E-09-7.86848040E-14    2
-4.05410765E+04-1.08505405E+02-2.95097578E+00+9.82464841E-02-7.59224537E-05    3
+2.92820284E-08-4.45657904E-12-3.08990846E+04+4.77269227E+01+0.00000000E+00    4
C6H11O13-2OOH           C   6H  12O   3    0G   300.000  5000.000 1425.000    51
+2.63085971E+01+2.61546948E-02-8.77769854E-06+1.34612150E-09-7.74534976E-14    2
-4.34234785E+04-1.10295283E+02-5.04452953E+00+1.05918270E-01-8.58242816E-05    3
+3.47733637E-08-5.55440543E-12-3.34375726E+04+5.53559272E+01+0.00000000E+00    4
C6H11O13-4OOH           C   6H  12O   3    0G   300.000  5000.000 1425.000    51
+2.63085971E+01+2.61546948E-02-8.77769854E-06+1.34612150E-09-7.74534976E-14    2
-4.34234785E+04-1.10295283E+02-5.04452953E+00+1.05918270E-01-8.58242816E-05    3
+3.47733637E-08-5.55440543E-12-3.34375726E+04+5.53559272E+01+0.00000000E+00    4
C6H11O13-5OOH           C   6H  12O   3    0G   300.000  5000.000 1425.000    51
+2.63085971E+01+2.61546948E-02-8.77769854E-06+1.34612150E-09-7.74534976E-14    2
-4.34234785E+04-1.10295283E+02-5.04452953E+00+1.05918270E-01-8.58242816E-05    3
+3.47733637E-08-5.55440543E-12-3.34375726E+04+5.53559272E+01+0.00000000E+00    4
C6H11O13-6OOH           C   6H  12O   3    0G   300.000  5000.000 1416.000    51
+2.54629106E+01+2.72623626E-02-9.24125642E-06+1.42660936E-09-8.24582230E-14    2
-4.12981961E+04-1.04829559E+02-5.60563964E+00+1.04991651E-01-8.32471205E-05    3
+3.31747712E-08-5.24343976E-12-3.12256985E+04+5.98605002E+01+0.00000000E+00    4
C6H11O14-2OOH           C   6H  12O   3    0G   300.000  5000.000 1425.000    41
+2.56382200E+01+2.71509666E-02-9.12183288E-06+1.39988818E-09-8.05862525E-14    2
-5.35027729E+04-1.08120825E+02-7.31154133E+00+1.11367218E-01-9.09451363E-05    3
+3.71421722E-08-5.98132077E-12-4.30436125E+04+6.58337228E+01+0.00000000E+00    4
C6H11O14-3OOH           C   6H  12O   3    0G   300.000  5000.000 1425.000    41
+2.56382200E+01+2.71509666E-02-9.12183288E-06+1.39988818E-09-8.05862525E-14    2
-5.35027729E+04-1.08120825E+02-7.31154133E+00+1.11367218E-01-9.09451363E-05    3
+3.71421722E-08-5.98132077E-12-4.30436125E+04+6.58337228E+01+0.00000000E+00    4
C6H11O14-5OOH           C   6H  12O   3    0G   300.000  5000.000 1425.000    41
+2.56382200E+01+2.71509666E-02-9.12183288E-06+1.39988818E-09-8.05862525E-14    2
-5.35027729E+04-1.08120825E+02-7.31154133E+00+1.11367218E-01-9.09451363E-05    3
+3.71421722E-08-5.98132077E-12-4.30436125E+04+6.58337228E+01+0.00000000E+00    4
C6H11O14-6OOH           C   6H  12O   3    0G   300.000  5000.000 1412.000    41
+2.45656595E+01+2.85283025E-02-9.69282356E-06+1.49844211E-09-8.66890301E-14    2
-5.12777917E+04-1.01359408E+02-9.39812599E+00+1.17516430E-01-9.95761400E-05    3
+4.27858226E-08-7.31024149E-12-4.06059311E+04+7.73575995E+01+0.00000000E+00    4
C6H11O15-2OOH           C   6H  12O   3    0G   300.000  5000.000 1413.000    31
+2.57514330E+01+2.79489406E-02-9.49498364E-06+1.46787433E-09-8.49251091E-14    2
-5.58563407E+04-1.13983278E+02-9.56356958E+00+1.21160691E-01-1.04208598E-04    3
+4.51613897E-08-7.75046859E-12-4.48492256E+04+7.15665603E+01+0.00000000E+00    4
C6H11O15-3OOH           C   6H  12O   3    0G   300.000  5000.000 1413.000    31
+2.57514330E+01+2.79489406E-02-9.49498364E-06+1.46787433E-09-8.49251091E-14    2
-5.58563407E+04-1.13983278E+02-9.56356958E+00+1.21160691E-01-1.04208598E-04    3
+4.51613897E-08-7.75046859E-12-4.48492256E+04+7.15665603E+01+0.00000000E+00    4
C6H11O15-4OOH           C   6H  12O   3    0G   300.000  5000.000 1413.000    31
+2.57514330E+01+2.79489406E-02-9.49498364E-06+1.46787433E-09-8.49251091E-14    2
-5.58563407E+04-1.13983278E+02-9.56356958E+00+1.21160691E-01-1.04208598E-04    3
+4.51613897E-08-7.75046859E-12-4.48492256E+04+7.15665603E+01+0.00000000E+00    4
C6H11O15-6OOH           C   6H  12O   3    0G   300.000  5000.000 1410.000    31
+2.50812660E+01+2.87541510E-02-9.82374389E-06+1.52441144E-09-8.84255093E-14    2
-5.37741881E+04-1.09448133E+02-9.86762792E+00+1.19225986E-01-1.00035576E-04    3
+4.24450450E-08-7.16631181E-12-4.26812046E+04+7.48455212E+01+0.00000000E+00    4
C6H11O23-1OOH           C   6H  12O   3    0G   300.000  5000.000 1425.000    61
+2.69564039E+01+2.52133315E-02-8.46015924E-06+1.29728465E-09-7.46387394E-14    2
-4.25735727E+04-1.11973745E+02-3.00051751E+00+1.01052251E-01-8.12852734E-05    3
+3.26822710E-08-5.17958864E-12-3.29962026E+04+4.64312180E+01+0.00000000E+00    4
C6H11O23-4OOH           C   6H  12O   3    0G   300.000  5000.000 1443.000    61
+2.80583928E+01+2.37928220E-02-7.87310190E-06+1.19630476E-09-6.84039421E-14    2
-4.48154981E+04-1.18929909E+02-2.32023655E+00+1.01282059E-01-8.24064664E-05    3
+3.31693978E-08-5.21408840E-12-3.52234339E+04+4.13949391E+01+0.00000000E+00    4
C6H11O23-5OOH           C   6H  12O   3    0G   300.000  5000.000 1443.000    61
+2.80583928E+01+2.37928220E-02-7.87310190E-06+1.19630476E-09-6.84039421E-14    2
-4.48154981E+04-1.18929909E+02-2.32023655E+00+1.01282059E-01-8.24064664E-05    3
+3.31693978E-08-5.21408840E-12-3.52234339E+04+4.13949391E+01+0.00000000E+00    4
C6H11O23-6OOH           C   6H  12O   3    0G   300.000  5000.000 1425.000    61
+2.69564039E+01+2.52133315E-02-8.46015924E-06+1.29728465E-09-7.46387394E-14    2
-4.25735727E+04-1.11973745E+02-3.00051751E+00+1.01052251E-01-8.12852734E-05    3
+3.26822710E-08-5.17958864E-12-3.29962026E+04+4.64312180E+01+0.00000000E+00    4
C6H11O24-1OOH           C   6H  12O   3    0G   300.000  5000.000 1423.000    51
+2.59111942E+01+2.64899573E-02-8.89134224E-06+1.36353586E-09-7.84507854E-14    2
-4.32925163E+04-1.07879889E+02-5.62254622E+00+1.07701280E-01-8.86273652E-05    3
+3.66476695E-08-5.99023124E-12-3.33282520E+04+5.84076967E+01+0.00000000E+00    4
C6H11O24-3OOH           C   6H  12O   3    0G   300.000  5000.000 1433.000    51
+2.68522312E+01+2.52818726E-02-8.39099827E-06+1.27724274E-09-7.31102872E-14    2
-4.54678687E+04-1.13918662E+02-5.05790795E+00+1.08518606E-01-9.08699191E-05    3
+3.79673868E-08-6.23050248E-12-3.55387589E+04+5.38980265E+01+0.00000000E+00    4
C6H11O24-5OOH           C   6H  12O   3    0G   300.000  5000.000 1433.000    51
+2.68522312E+01+2.52818726E-02-8.39099827E-06+1.27724274E-09-7.31102872E-14    2
-4.54678687E+04-1.13918662E+02-5.05790795E+00+1.08518606E-01-9.08699191E-05    3
+3.79673868E-08-6.23050248E-12-3.55387589E+04+5.38980265E+01+0.00000000E+00    4
C6H11O24-6OOH           C   6H  12O   3    0G   300.000  5000.000 1423.000    51
+2.59111942E+01+2.64899573E-02-8.89134224E-06+1.36353586E-09-7.84507854E-14    2
-4.32925163E+04-1.07879889E+02-5.62254622E+00+1.07701280E-01-8.86273652E-05    3
+3.66476695E-08-5.99023124E-12-3.33282520E+04+5.84076967E+01+0.00000000E+00    4
C6H11O25-1OOH           C   6H  12O   3    0G   300.000  5000.000 1416.000    41
+2.48755287E+01+2.78565097E-02-9.37289923E-06+1.43948573E-09-8.28962898E-14    2
-5.32048100E+04-1.03584543E+02-9.24035424E+00+1.19425795E-01-1.03974569E-04    3
+4.57446356E-08-7.95660813E-12-4.27327015E+04+7.51088527E+01+0.00000000E+00    4
C6H11O25-3OOH           C   6H  12O   3    0G   300.000  5000.000 1421.000    41
+2.54725769E+01+2.68960204E-02-8.94476389E-06+1.36283531E-09-7.80436306E-14    2
-5.51746673E+04-1.07502255E+02-8.92888836E+00+1.22020603E-01-1.09968258E-04    3
+4.98119645E-08-8.85746002E-12-4.49187054E+04+7.16554572E+01+0.00000000E+00    4
C6H11O34-1OOH           C   6H  12O   3    0G   300.000  5000.000 1425.000    61
+2.69564039E+01+2.52133315E-02-8.46015924E-06+1.29728465E-09-7.46387394E-14    2
-4.25735727E+04-1.11973745E+02-3.00051751E+00+1.01052251E-01-8.12852734E-05    3
+3.26822710E-08-5.17958864E-12-3.29962026E+04+4.64312180E+01+0.00000000E+00    4
C6H11O34-2OOH           C   6H  12O   3    0G   300.000  5000.000 1443.000    61
+2.80583928E+01+2.37928220E-02-7.87310190E-06+1.19630476E-09-6.84039421E-14    2
-4.48154981E+04-1.18929909E+02-2.32023655E+00+1.01282059E-01-8.24064664E-05    3
+3.31693978E-08-5.21408840E-12-3.52234339E+04+4.13949391E+01+0.00000000E+00    4
C5H9O12-5               C   5H   9O   1    0G   300.000  5000.000 1428.000    31
+1.71692866E+01+1.96439921E-02-6.56270756E-06+1.00313537E-09-5.75797826E-14    2
+1.20372734E+02-6.41594420E+01-4.74570948E+00+7.55874963E-02-6.08534529E-05    3
+2.46895048E-08-3.96232760E-12+7.08653513E+03+5.15668737E+01+0.00000000E+00    4
C4H7O12-4               C   4H   7O   1    0G   300.000  5000.000 1521.000    21
+1.34570917E+01+1.40456552E-02-4.31981858E-06+6.22563489E-10-3.42463069E-14    2
+4.88696367E+03-4.44520295E+01-3.37974855E+00+6.03280881E-02-5.19900485E-05    3
+2.23629697E-08-3.72920327E-12+9.80004298E+03+4.31033481E+01+0.00000000E+00    4
C4H7O13-4               C   4H   7O   1    0G   300.000  5000.000 1436.000    11
+1.26383103E+01+1.59453761E-02-5.13309123E-06+7.64898728E-10-4.31253622E-14    2
+3.91648984E+03-4.20740863E+01-4.66267157E+00+6.15207910E-02-5.06948989E-05    3
+2.11863240E-08-3.49163560E-12+9.24461326E+03+4.87364061E+01+0.00000000E+00    4
C4H7O23-1               C   4H   7O   1    0G   300.000  5000.000 1324.000    21
+8.53917898E+00+1.94224428E-02-6.06403336E-06+6.79865833E-10-1.50192364E-14    2
+5.95005552E+03-1.55618089E+01-3.45625302E+00+6.17954277E-02-5.36422388E-05    3
+2.24943234E-08-3.70306875E-12+7.74377568E+03+4.22227921E+01+0.00000000E+00    4
C5H9O13-5               C   5H   9O   1    0G   300.000  5000.000 1458.000    21
+1.55990028E+01+2.00371413E-02-6.41154602E-06+9.50807571E-10-5.34042125E-14    2
+3.37602077E+00-5.60383294E+01-6.25393631E+00+7.92184870E-02-6.70994450E-05    3
+2.87608390E-08-4.83752138E-12+6.54668516E+03+5.80476602E+01+0.00000000E+00    4
C5H9O14-5               C   5H   9O   1    0G   300.000  5000.000 1447.000    11
+1.54610559E+01+2.06809909E-02-6.66141956E-06+9.93099401E-10-5.60118090E-14    2
-1.03327057E+04-5.70023035E+01-7.49219030E+00+8.07085780E-02-6.60336535E-05    3
+2.72423613E-08-4.41750289E-12-3.23749643E+03+6.36020351E+01+0.00000000E+00    4
C5H9O23-1               C   5H   9O   1    0G   300.000  5000.000 1424.000    31
+1.77401551E+01+1.92298085E-02-6.43473125E-06+9.84654362E-10-5.65624830E-14    2
-2.05448135E+03-6.82408862E+01-4.67636252E+00+7.74809264E-02-6.42244373E-05    3
+2.68440080E-08-4.43868315E-12+4.97926865E+03+4.97877901E+01+0.00000000E+00    4
C5H9O23-5               C   5H   9O   1    0G   300.000  5000.000 1424.000    31
+1.77401551E+01+1.92298085E-02-6.43473125E-06+9.84654362E-10-5.65624830E-14    2
-2.05448135E+03-6.82408862E+01-4.67636252E+00+7.74809264E-02-6.42244373E-05    3
+2.68440080E-08-4.43868315E-12+4.97926865E+03+4.97877901E+01+0.00000000E+00    4
C5H9O24-1               C   5H   9O   1    0G   300.000  5000.000 1398.000    21
+1.40157807E+01+2.51554423E-02-1.11149003E-05+2.14885206E-09-1.44559627E-13    2
-1.54769089E+03-4.88521063E+01-6.45048964E+00+8.25684509E-02-7.30635550E-05    3
+3.23767886E-08-5.72480023E-12+4.47417427E+03+5.74524602E+01+0.00000000E+00    4
C6KET12O                C   6H  11O   2    0G   300.000  5000.000 1380.000    51
+2.44011335E+01+2.43695802E-02-8.52760748E-06+1.34452656E-09-7.88560069E-14    2
-3.46915506E+04-9.76141351E+01+2.48709886E+00+6.84851704E-02-3.91082619E-05    3
+9.26081053E-09-5.01384589E-13-2.64222925E+04+2.25084325E+01+0.00000000E+00    4
C6KET13O                C   6H  11O   2    0G   300.000  5000.000 1420.000    51
+2.43086453E+01+2.35169486E-02-8.03437802E-06+1.24733142E-09-7.23954247E-14    2
-3.52041500E+04-9.76594163E+01+3.39465791E+00+6.34450550E-02-3.11900396E-05    3
+3.70312592E-09+8.80779018E-13-2.72582338E+04+1.74777979E+01+0.00000000E+00    4
C6KET14O                C   6H  11O   2    0G   300.000  5000.000 1420.000    51
+2.43086453E+01+2.35169486E-02-8.03437802E-06+1.24733142E-09-7.23954247E-14    2
-3.52041500E+04-9.76594163E+01+3.39465791E+00+6.34450550E-02-3.11900396E-05    3
+3.70312592E-09+8.80779018E-13-2.72582338E+04+1.74777979E+01+0.00000000E+00    4
C6KET15O                C   6H  11O   2    0G   300.000  5000.000 1420.000    51
+2.43086453E+01+2.35169486E-02-8.03437802E-06+1.24733142E-09-7.23954247E-14    2
-3.52041500E+04-9.76594163E+01+3.39465791E+00+6.34450550E-02-3.11900396E-05    3
+3.70312592E-09+8.80779018E-13-2.72582338E+04+1.74777979E+01+0.00000000E+00    4
C6KET21O                C   6H  11O   2    0G   300.000  5000.000 1487.000    51
+2.25293622E+01+2.47975925E-02-8.43579282E-06+1.30658010E-09-7.57309929E-14    2
-3.53514289E+04-8.65954633E+01+7.39116829E+00+4.44580281E-02-6.38228035E-06    3
-9.61459324E-09+3.45678863E-12-2.86152512E+04+1.28093150E-01+0.00000000E+00    4
C6KET23O                C   6H  11O   2    0G   300.000  5000.000 1386.000    51
+2.29408073E+01+2.51899756E-02-8.71525786E-06+1.36369341E-09-7.95562705E-14    2
-3.77254587E+04-8.90236293E+01+3.25181786E+00+6.46413698E-02-3.58852109E-05    3
+8.30469730E-09-4.25746250E-13-3.02655065E+04+1.89862996E+01+0.00000000E+00    4
C6KET24O                C   6H  11O   2    0G   300.000  5000.000 1530.000    51
+2.17184075E+01+2.47007497E-02-8.21787847E-06+1.25253279E-09-7.17484997E-14    2
-3.75473266E+04-8.19767338E+01+4.41342175E+00+5.98412718E-02-3.19612065E-05    3
+6.55909263E-09-5.07843738E-14-3.11596284E+04+1.25825004E+01+0.00000000E+00    4
C6KET25O                C   6H  11O   2    0G   300.000  5000.000 1530.000    51
+2.17184075E+01+2.47007497E-02-8.21787847E-06+1.25253279E-09-7.17484997E-14    2
-3.75473266E+04-8.19767338E+01+4.41342175E+00+5.98412718E-02-3.19612065E-05    3
+6.55909263E-09-5.07843738E-14-3.11596284E+04+1.25825004E+01+0.00000000E+00    4
C6KET26O                C   6H  11O   2    0G   300.000  5000.000 1527.000    51
+2.13007803E+01+2.58716731E-02-8.79653453E-06+1.36062148E-09-7.87479444E-14    2
-3.57843109E+04-7.96089891E+01+4.01263738E+00+5.66756784E-02-2.38571625E-05    3
+8.77122160E-10+1.22542395E-12-2.89322231E+04+1.64535234E+01+0.00000000E+00    4
C6KET31O                C   6H  11O   2    0G   300.000  5000.000 1305.000    51
+2.20864552E+01+2.46779992E-02-8.28346973E-06+1.27113585E-09-7.31921565E-14    2
-3.61540517E+04-8.46188998E+01+5.02858055E+00+5.12156892E-02-1.40537055E-05    3
-6.12620240E-09+2.92422949E-12-2.91213820E+04+1.13420391E+01+0.00000000E+00    4
C6KET32O                C   6H  11O   2    0G   300.000  5000.000 1381.000    51
+2.23075626E+01+2.54572934E-02-8.74888878E-06+1.36294097E-09-7.92726719E-14    2
-3.75305099E+04-8.59089550E+01+4.28777527E+00+5.83079361E-02-2.63826419E-05    3
+2.44071634E-09+8.67814900E-13-3.04212126E+04+1.40253081E+01+0.00000000E+00    4
C6KET34O                C   6H  11O   2    0G   300.000  5000.000 1381.000    51
+2.23075626E+01+2.54572934E-02-8.74888878E-06+1.36294097E-09-7.92726719E-14    2
-3.75305099E+04-8.59089550E+01+4.28777527E+00+5.83079361E-02-2.63826419E-05    3
+2.44071634E-09+8.67814900E-13-3.04212126E+04+1.40253081E+01+0.00000000E+00    4
C6KET35O                C   6H  11O   2    0G   300.000  5000.000 1416.000    51
+2.26318948E+01+2.41684263E-02-8.10341688E-06+1.24303233E-09-7.15692685E-14    2
-3.84096424E+04-8.87241802E+01+4.84610323E+00+5.24943003E-02-1.55391890E-05    3
-5.44987122E-09+2.81073621E-12-3.11401488E+04+1.11045620E+01+0.00000000E+00    4
C6KET36O                C   6H  11O   2    0G   300.000  5000.000 1305.000    51
+2.20864552E+01+2.46779992E-02-8.28346973E-06+1.27113585E-09-7.31921565E-14    2
-3.61540517E+04-8.46188998E+01+5.02858055E+00+5.12156892E-02-1.40537055E-05    3
-6.12620240E-09+2.92422949E-12-2.91213820E+04+1.13420391E+01+0.00000000E+00    4
C6H12OOH1-2O            C   6H  13O   3    0G   300.000  5000.000 1535.000    71
+2.92647989E+01+2.69146554E-02-9.38475487E-06+1.47659709E-09-8.64902012E-14    2
-3.71424073E+04-1.22240832E+02+2.80591255E+00+7.79229941E-02-4.02499146E-05    3
+6.01126951E-09+7.21748984E-13-2.70819447E+04+2.33451434E+01+0.00000000E+00    4
C6H12OOH1-3O            C   6H  13O   3    0G   300.000  5000.000 1535.000    71
+2.92647989E+01+2.69146554E-02-9.38475487E-06+1.47659709E-09-8.64902012E-14    2
-3.71424073E+04-1.22240832E+02+2.80591255E+00+7.79229941E-02-4.02499146E-05    3
+6.01126951E-09+7.21748984E-13-2.70819447E+04+2.33451434E+01+0.00000000E+00    4
C6H12OOH1-4O            C   6H  13O   3    0G   300.000  5000.000 1535.000    71
+2.92647989E+01+2.69146554E-02-9.38475487E-06+1.47659709E-09-8.64902012E-14    2
-3.71424073E+04-1.22240832E+02+2.80591255E+00+7.79229941E-02-4.02499146E-05    3
+6.01126951E-09+7.21748984E-13-2.70819447E+04+2.33451434E+01+0.00000000E+00    4
C6H12OOH1-5O            C   6H  13O   3    0G   300.000  5000.000 1535.000    71
+2.92647989E+01+2.69146554E-02-9.38475487E-06+1.47659709E-09-8.64902012E-14    2
-3.71424073E+04-1.22240832E+02+2.80591255E+00+7.79229941E-02-4.02499146E-05    3
+6.01126951E-09+7.21748984E-13-2.70819447E+04+2.33451434E+01+0.00000000E+00    4
C6H12OOH2-1O            C   6H  13O   3    0G   300.000  5000.000 1409.000    71
+2.68394200E+01+2.78771803E-02-9.46581223E-06+1.46245818E-09-8.45621758E-14    2
-3.54171892E+04-1.06763190E+02+3.34629056E+00+8.24137185E-02-5.70430278E-05    3
+1.99491279E-08-2.77573029E-12-2.73151509E+04+1.93763739E+01+0.00000000E+00    4
C6H12OOH2-3O            C   6H  13O   3    0G   300.000  5000.000 1408.000    71
+2.70100981E+01+2.75803123E-02-9.32839137E-06+1.43724826E-09-8.29386001E-14    2
-3.73322411E+04-1.08327965E+02+2.14026689E+00+9.05994482E-02-7.11844189E-05    3
+2.92349633E-08-4.87305224E-12-2.92400104E+04+2.34016654E+01+0.00000000E+00    4
C6H12OOH2-4O            C   6H  13O   3    0G   300.000  5000.000 1408.000    71
+2.70100981E+01+2.75803123E-02-9.32839137E-06+1.43724826E-09-8.29386001E-14    2
-3.73322411E+04-1.08327965E+02+2.14026689E+00+9.05994482E-02-7.11844189E-05    3
+2.92349633E-08-4.87305224E-12-2.92400104E+04+2.34016654E+01+0.00000000E+00    4
C6H12OOH2-5O            C   6H  13O   3    0G   300.000  5000.000 1408.000    71
+2.70100981E+01+2.75803123E-02-9.32839137E-06+1.43724826E-09-8.29386001E-14    2
-3.73322411E+04-1.08327965E+02+2.14026689E+00+9.05994482E-02-7.11844189E-05    3
+2.92349633E-08-4.87305224E-12-2.92400104E+04+2.34016654E+01+0.00000000E+00    4
C6H12OOH2-6O            C   6H  13O   3    0G   300.000  5000.000 1409.000    71
+2.68394200E+01+2.78771803E-02-9.46581223E-06+1.46245818E-09-8.45621758E-14    2
-3.54171892E+04-1.06763190E+02+3.34629056E+00+8.24137185E-02-5.70430278E-05    3
+1.99491279E-08-2.77573029E-12-2.73151509E+04+1.93763739E+01+0.00000000E+00    4
C6H12OOH3-1O            C   6H  13O   3    0G   300.000  5000.000 1409.000    71
+2.68394200E+01+2.78771803E-02-9.46581223E-06+1.46245818E-09-8.45621758E-14    2
-3.54171892E+04-1.06763190E+02+3.34629056E+00+8.24137185E-02-5.70430278E-05    3
+1.99491279E-08-2.77573029E-12-2.73151509E+04+1.93763739E+01+0.00000000E+00    4
C6H12OOH3-2O            C   6H  13O   3    0G   300.000  5000.000 1408.000    71
+2.70100981E+01+2.75803123E-02-9.32839137E-06+1.43724826E-09-8.29386001E-14    2
-3.73322411E+04-1.08327965E+02+2.14026689E+00+9.05994482E-02-7.11844189E-05    3
+2.92349633E-08-4.87305224E-12-2.92400104E+04+2.34016654E+01+0.00000000E+00    4
C6H12OOH3-4O            C   6H  13O   3    0G   300.000  5000.000 1408.000    71
+2.70100981E+01+2.75803123E-02-9.32839137E-06+1.43724826E-09-8.29386001E-14    2
-3.73322411E+04-1.08327965E+02+2.14026689E+00+9.05994482E-02-7.11844189E-05    3
+2.92349633E-08-4.87305224E-12-2.92400104E+04+2.34016654E+01+0.00000000E+00    4
C6H12OOH3-5O            C   6H  13O   3    0G   300.000  5000.000 1408.000    71
+2.70100981E+01+2.75803123E-02-9.32839137E-06+1.43724826E-09-8.29386001E-14    2
-3.73322411E+04-1.08327965E+02+2.14026689E+00+9.05994482E-02-7.11844189E-05    3
+2.92349633E-08-4.87305224E-12-2.92400104E+04+2.34016654E+01+0.00000000E+00    4
C6H12OOH3-6O            C   6H  13O   3    0G   300.000  5000.000 1409.000    71
+2.68394200E+01+2.78771803E-02-9.46581223E-06+1.46245818E-09-8.45621758E-14    2
-3.54171892E+04-1.06763190E+02+3.34629056E+00+8.24137185E-02-5.70430278E-05    3
+1.99491279E-08-2.77573029E-12-2.73151509E+04+1.93763739E+01+0.00000000E+00    4
C6Y2                    C   6H  12O   1    0G   300.000  5000.000 1393.000    51
+1.91702580E+01+2.71941021E-02-9.14602800E-06+1.40414058E-09-8.08375794E-14    2
-4.34193894E+04-7.21956796E+01+1.91874702E+00+6.12265198E-02-3.15172753E-05    3
+6.28658563E-09-6.56228984E-14-3.68622671E+04+2.25762120E+01+0.00000000E+00    4
CH3COOH           G 6/00C  2.H  4.O  2.   0.G   200.000  6000.000 1000.        1
+7.67084601E+00+1.35152602E-02-5.25874333E-06+8.93184479E-10-5.53180543E-14    2
-5.57560970E+04-1.54677315E+01+2.78950201E+00+9.99941719E-03+3.42572245E-05    3
-5.09031329E-08+2.06222185E-11-5.34752488E+04+1.41053123E+01-5.19873137E+04    4
C2H5COOH          T11/07C  3.H  6.O  2.   0.G   200.000  6000.000 1000.        1
+8.61036813E+00+1.87894582E-02-6.70711294E-06+1.07428300E-09-6.38870386E-14    2
-5.84807549E+04-1.63110488E+01+5.51515351E+00-1.02654246E-05+7.54897239E-05    3
-9.81744541E-08+3.88829515E-11-5.63618075E+04+6.11744431E+00-5.42266279E+04    4
C6H12-1                 C   6H  12    0    0G   300.000  5000.000 1391.000    41
+1.77068656E+01+2.69421757E-02-9.19125439E-06+1.42442840E-09-8.25377749E-14    2
-1.41883983E+04-6.77121636E+01-4.88101166E-01+6.60223990E-02-4.03430121E-05    3
+1.23616901E-08-1.50560345E-12-7.49399629E+03+3.12755041E+01+0.00000000E+00    4
C6H12-2                 C   6H  12    0    0G   300.000  5000.000 1388.000    41
+1.72811801E+01+2.72154214E-02-9.26717645E-06+1.43446313E-09-8.30514585E-14    2
-1.53826845E+04-6.59650838E+01+2.64795074E-01+6.14938008E-02-3.36108501E-05    3
+8.31993597E-09-6.42021164E-13-8.89772499E+03+2.74114997E+01+0.00000000E+00    4
C6H12-3                 C   6H  12    0    0G   300.000  5000.000 1386.000    41
+1.70313735E+01+2.73270171E-02-9.28504971E-06+1.43523149E-09-8.30182955E-14    2
-1.53031077E+04-6.53708588E+01-1.72607040E-01+6.19357715E-02-3.37261047E-05    3
+8.23624938E-09-6.03434172E-13-8.75056335E+03+2.90378440E+01+0.00000000E+00    4
C6H111-3                C   6H  11    0    0G   300.000  5000.000 1380.000    31
+1.81062746E+01+2.41474871E-02-8.16683437E-06+1.25923677E-09-7.27359868E-14    2
+2.45878515E+03-6.97527464E+01-1.80747803E-01+6.22067565E-02-3.63722507E-05    3
+9.77864452E-09-8.75066308E-13+9.24216018E+03+3.00591380E+01+0.00000000E+00    4
C6H111-4                C   6H  11    0    0G   300.000  5000.000 1393.000    41
+1.61989292E+01+2.55342673E-02-8.67483385E-06+1.34064100E-09-7.75312952E-14    2
+9.67127430E+03-5.61196642E+01+1.15589239E+00+5.34977768E-02-2.48120970E-05    3
+3.38660024E-09+4.19889741E-13+1.55875202E+04+2.71720322E+01+0.00000000E+00    4
C6H111-5                C   6H  11    0    0G   300.000  5000.000 1393.000    41
+1.61989292E+01+2.55342673E-02-8.67483385E-06+1.34064100E-09-7.75312952E-14    2
+9.67127430E+03-5.61196642E+01+1.15589239E+00+5.34977768E-02-2.48120970E-05    3
+3.38660024E-09+4.19889741E-13+1.55875202E+04+2.71720322E+01+0.00000000E+00    4
C6H111-6                C   6H  11    0    0G   300.000  5000.000 1387.000    51
+1.74644753E+01+2.47005987E-02-8.53334148E-06+1.33367297E-09-7.77343118E-14    2
+1.07088778E+04-6.39032857E+01+8.71879475E-02+6.14727795E-02-3.75054886E-05    3
+1.14767733E-08-1.41643272E-12+1.71987905E+04+3.09015588E+01+0.00000000E+00    4
C6H112-4                C   6H  11    0    0G   300.000  5000.000 1388.000    31
+1.68906239E+01+2.55067554E-02-8.69671971E-06+1.34743880E-09-7.80675027E-14    2
+1.66448555E+03-6.50840113E+01-8.09214028E-02+6.00167919E-02-3.34681107E-05    3
+8.44580243E-09-6.67121954E-13+8.07876099E+03+2.78967527E+01+0.00000000E+00    4
C6H112-5                C   6H  11    0    0G   300.000  5000.000 1385.000    41
+1.57816863E+01+2.57956633E-02-8.74566769E-06+1.34977950E-09-7.79887258E-14    2
+8.48313934E+03-5.43988313E+01+2.08038945E+00+4.83569471E-02-1.72566989E-05    3
-1.13784525E-09+1.38654068E-12+1.41534725E+04+2.24803229E+01+0.00000000E+00    4
C6H112-6                C   6H  11    0    0G   300.000  5000.000 1385.000    51
+1.69591869E+01+2.51413831E-02-8.68761395E-06+1.35795747E-09-7.91556719E-14    2
+9.53673982E+03-6.17306897E+01+6.38205633E-01+5.78758020E-02-3.22194721E-05    3
+8.38982851E-09-7.74542374E-13+1.58248386E+04+2.79713260E+01+0.00000000E+00    4
C6H113-1                C   6H  11    0    0G   300.000  5000.000 1387.000    41
+1.63801476E+01+2.54479755E-02-8.66105290E-06+1.34023418E-09-7.75806403E-14    2
+9.84382560E+03-5.83757912E+01+2.39410938E-01+5.82991009E-02-3.24715921E-05    3
+8.38108128E-09-7.27332655E-13+1.59623764E+04+3.00781535E+01+0.00000000E+00    4
C6H12OH-1J2             C   6H  13O   1    0G   300.000  5000.000 1395.000    61
+2.05219095E+01+2.85941986E-02-9.71574333E-06+1.50154769E-09-8.68352394E-14    2
-2.46176531E+04-7.58039610E+01+1.52879690E+00+7.02411418E-02-4.39606425E-05    3
+1.40750120E-08-1.82860462E-12-1.77206486E+04+2.72130211E+01+0.00000000E+00    4
C6H12OH-2J1             C   6H  13O   1    0G   300.000  5000.000 1403.000    61
+2.16778753E+01+2.71851643E-02-9.13650238E-06+1.40152530E-09-8.06255019E-14    2
-2.55354913E+04-8.29034809E+01+1.12882665E+00+7.79334290E-02-5.78628264E-05    3
+2.29540709E-08-3.76055142E-12-1.86725358E+04+2.64835374E+01+0.00000000E+00    4
C6H12OH-2J3             C   6H  13O   1    0G   300.000  5000.000 1402.000    61
+2.08484871E+01+2.76635202E-02-9.25462670E-06+1.41532103E-09-8.12482889E-14    2
-2.65002333E+04-7.79996791E+01+1.24040698E+00+7.41986609E-02-5.16292083E-05    3
+1.90231170E-08-2.89350308E-12-1.97802722E+04+2.70192329E+01+0.00000000E+00    4
C6H12OH-3J2             C   6H  13O   1    0G   300.000  5000.000 1402.000    61
+2.08484871E+01+2.76635202E-02-9.25462670E-06+1.41532103E-09-8.12482889E-14    2
-2.65002333E+04-7.79996791E+01+1.24040698E+00+7.41986609E-02-5.16292083E-05    3
+1.90231170E-08-2.89350308E-12-1.97802722E+04+2.70192329E+01+0.00000000E+00    4
C6H12OH-3J4             C   6H  13O   1    0G   300.000  5000.000 1402.000    61
+2.08484871E+01+2.76635202E-02-9.25462670E-06+1.41532103E-09-8.12482889E-14    2
-2.65002333E+04-7.79996791E+01+1.24040698E+00+7.41986609E-02-5.16292083E-05    3
+1.90231170E-08-2.89350308E-12-1.97802722E+04+2.70192329E+01+0.00000000E+00    4
C6H12OH-1O2-2           C   6H  13O   3    0G   300.000  5000.000 1404.000    71
+2.62416220E+01+2.83873841E-02-9.64269140E-06+1.49018659E-09-8.61823559E-14    2
-4.52283711E+04-1.03056223E+02+1.21185034E+00+8.86935209E-02-6.52629776E-05    3
+2.48084263E-08-3.82705801E-12-3.67836493E+04+3.06087511E+01+0.00000000E+00    4
C6H12OH-2O2-1           C   6H  13O   3    0G   300.000  5000.000 1402.000    71
+2.54686767E+01+2.90602674E-02-9.87649038E-06+1.52670395E-09-8.83047932E-14    2
-4.49414723E+04-9.84561539E+01+8.48833477E-01+8.96057240E-02-6.76377691E-05    3
+2.68760659E-08-4.38117112E-12-3.67038364E+04+3.26746588E+01+0.00000000E+00    4
C6H12OH-2O2-3           C   6H  13O   3    0G   300.000  5000.000 1409.000    71
+2.58464390E+01+2.81918402E-02-9.45730022E-06+1.44892549E-09-8.32798272E-14    2
-4.67848660E+04-1.01026245E+02+1.25084224E+00+9.16687695E-02-7.30413883E-05    3
+3.06072325E-08-5.20205053E-12-3.88977871E+04+2.88405166E+01+0.00000000E+00    4
C6H12OH-3O2-2           C   6H  13O   3    0G   300.000  5000.000 1409.000    71
+2.58464390E+01+2.81918402E-02-9.45730022E-06+1.44892549E-09-8.32798272E-14    2
-4.67848660E+04-1.01026245E+02+1.25084224E+00+9.16687695E-02-7.30413883E-05    3
+3.06072325E-08-5.20205053E-12-3.88977871E+04+2.88405166E+01+0.00000000E+00    4
C6H12OH-3O2-4           C   6H  13O   3    0G   300.000  5000.000 1409.000    71
+2.58464390E+01+2.81918402E-02-9.45730022E-06+1.44892549E-09-8.32798272E-14    2
-4.67848660E+04-1.01026245E+02+1.25084224E+00+9.16687695E-02-7.30413883E-05    3
+3.06072325E-08-5.20205053E-12-3.88977871E+04+2.88405166E+01+0.00000000E+00    4
C6H11-1D3O              C   6H  11O   1    0G   300.000  5000.000 1383.000    41
+2.12331424E+01+2.48369812E-02-8.66311197E-06+1.36270774E-09-7.97852110E-14    2
-8.51940477E+03-8.30721992E+01+2.10835922E+00+6.53603616E-02-4.08332113E-05    3
+1.28408111E-08-1.65145256E-12-1.36559988E+03+2.12769181E+01+0.00000000E+00    4
C6H11-1D4O              C   6H  11O   1    0G   300.000  5000.000 1407.000    41
+2.02215422E+01+2.43935819E-02-8.22353442E-06+1.26435910E-09-7.28591420E-14    2
-8.25970727E+03-7.72129963E+01+1.74896641E+00+6.59595125E-02-4.28715185E-05    3
+1.38805462E-08-1.74690339E-12-1.75725189E+03+2.24374197E+01+0.00000000E+00    4
C6H11-1D5O              C   6H  11O   1    0G   300.000  5000.000 1407.000    41
+2.02215422E+01+2.43935819E-02-8.22353442E-06+1.26435910E-09-7.28591420E-14    2
-8.25970727E+03-7.72129963E+01+1.74896641E+00+6.59595125E-02-4.28715185E-05    3
+1.38805462E-08-1.74690339E-12-1.75725189E+03+2.24374197E+01+0.00000000E+00    4
C6H11-1D6O              C   6H  11O   1    0G   300.000  5000.000 1394.000    41
+2.04129591E+01+2.48384017E-02-8.51026795E-06+1.32292012E-09-7.68252415E-14    2
-6.61087614E+03-7.80582419E+01+1.65674953E+00+6.36239531E-02-3.67332362E-05    3
+9.43984310E-09-7.26849847E-13+3.56296910E+02+2.43747538E+01+0.00000000E+00    4
C6H11-2D1O              C   6H  11O   1    0G   300.000  5000.000 1999.000    41
+1.63147059E+01+3.08756722E-02-1.12659286E-05+1.83193378E-09-1.09891277E-13    2
-5.48521972E+03-5.49439851E+01+6.40521825E+00+4.23558507E-02-7.63213993E-06    3
-5.93172496E-09+2.04790110E-12-1.07194029E+03+2.22105053E+00+0.00000000E+00    4
C6H11-2D4O              C   6H  11O   1    0G   300.000  5000.000 1380.000    41
+2.07337615E+01+2.52406898E-02-8.79759458E-06+1.38318161E-09-8.09557361E-14    2
-9.67476730E+03-8.08901300E+01+2.99930917E+00+6.04876255E-02-3.38261990E-05    3
+8.74283850E-09-7.93336016E-13-2.79750804E+03+1.67172352E+01+0.00000000E+00    4
C6H11-2D5O              C   6H  11O   1    0G   300.000  5000.000 1403.000    41
+1.98339795E+01+2.46335527E-02-8.28848420E-06+1.27278690E-09-7.32851452E-14    2
-9.47274334E+03-7.56901783E+01+2.54000411E+00+6.12908043E-02-3.59176813E-05    3
+9.70008242E-09-8.53771601E-13-3.16782333E+03+1.83891887E+01+0.00000000E+00    4
C6H11-2D6O              C   6H  11O   1    0G   300.000  5000.000 1390.000    41
+1.95292766E+01+2.55039957E-02-8.72047811E-06+1.35366557E-09-7.85302933E-14    2
-7.59824209E+03-7.36136387E+01+2.70082133E+00+5.78441974E-02-2.89980180E-05    3
+5.19918235E-09+1.16017596E-13-1.08709477E+03+1.91870295E+01+0.00000000E+00    4
C6H11-3D1O              C   6H  11O   1    0G   300.000  5000.000 1387.000    41
+1.92747614E+01+2.56242111E-02-8.74228366E-06+1.35514342E-09-7.85422000E-14    2
-7.51901058E+03-7.23056917E+01+2.34238003E+00+5.79452100E-02-2.86377646E-05    3
+4.84570137E-09+2.08901971E-13-9.52014318E+02+2.11357667E+01+0.00000000E+00    4
C6H11-3D2O              C   6H  11O   1    0G   300.000  5000.000 1380.000    41
+2.03827442E+01+2.55217123E-02-8.89072063E-06+1.39731901E-09-8.17627196E-14    2
-9.57080422E+03-7.90711932E+01+2.54762399E+00+6.07926451E-02-3.36415232E-05    3
+8.47505102E-09-7.17131188E-13-2.64230465E+03+1.91434934E+01+0.00000000E+00    4
NC5H11CHO               C   6H  12O   1    0G   300.000  5000.000 1387.000    51
+2.04873253E+01+2.68430457E-02-9.19116692E-06+1.42823241E-09-8.29221047E-14    2
-4.03782423E+04-8.01141801E+01+1.26510376E+00+6.45800926E-02-3.38952057E-05    3
+6.81908963E-09-7.71461981E-14-3.30370410E+04+2.55776945E+01+0.00000000E+00    4
NC5H11CO                C   6H  11O   1    0G   300.000  5000.000 1387.000    51
+2.00712533E+01+2.47109029E-02-8.46937882E-06+1.31698154E-09-7.65012214E-14    2
-2.14161547E+04-7.62093348E+01+2.03899694E+00+5.97834497E-02-3.08487256E-05    3
+5.75699235E-09+8.35477271E-14-1.45087642E+04+2.30358058E+01+0.00000000E+00    4
NC5H10CHO-1             C   6H  11O   1    0G   300.000  5000.000 1393.000    51
+2.06482100E+01+2.43700759E-02-8.38484086E-06+1.30722981E-09-7.60729502E-14    2
-2.02725848E+04-8.15155501E+01+5.78184620E-01+6.55176768E-02-3.75505403E-05    3
+9.10037088E-09-5.32652119E-13-1.28157111E+04+2.81624025E+01+0.00000000E+00    4
NC5H10CHO-2             C   6H  11O   1    0G   300.000  5000.000 1372.000    51
+1.91787632E+01+2.51424561E-02-8.54947751E-06+1.32258961E-09-7.65569904E-14    2
-1.65995988E+04-6.96557486E+01+2.74720823E+00+5.26109114E-02-1.88709415E-05    3
-2.03156157E-09+1.85276474E-12-9.92771663E+03+2.22524075E+01+0.00000000E+00    4
NC5H10CHO-3             C   6H  11O   1    0G   300.000  5000.000 1372.000    51
+1.91787632E+01+2.51424561E-02-8.54947751E-06+1.32258961E-09-7.65569904E-14    2
-1.65995988E+04-6.96557486E+01+2.74720823E+00+5.26109114E-02-1.88709415E-05    3
-2.03156157E-09+1.85276474E-12-9.92771663E+03+2.22524075E+01+0.00000000E+00    4
NC5H10CHO-4             C   6H  11O   1    0G   300.000  5000.000 1372.000    51
+1.91787632E+01+2.51424561E-02-8.54947751E-06+1.32258961E-09-7.65569904E-14    2
-1.65995988E+04-6.96557486E+01+2.74720823E+00+5.26109114E-02-1.88709415E-05    3
-2.03156157E-09+1.85276474E-12-9.92771663E+03+2.22524075E+01+0.00000000E+00    4
NC5H10CHO-5             C   6H  11O   1    0G   300.000  5000.000 1388.000    51
+1.99255677E+01+2.47873156E-02-8.48543707E-06+1.31842819E-09-7.65429548E-14    2
-1.52547493E+04-7.42913571E+01+1.60690963E+00+6.12092931E-02-3.29226741E-05    3
+7.03661827E-09-1.96773498E-13-8.31263906E+03+2.62561430E+01+0.00000000E+00    4
C6H10D13                C   6H  10    0    0G   300.000  5000.000 1395.000    31
+1.69088929E+01+2.30881104E-02-7.89077821E-06+1.22430123E-09-7.09963130E-14    2
-1.64475595E+03-6.46806187E+01-1.48701712E+00+6.83526916E-02-5.17682192E-05    3
+2.10789514E-08-3.57266133E-12+4.58162436E+03+3.34156371E+01+0.00000000E+00    4
C6H10D24                C   6H  10    0    0G   300.000  5000.000 1393.000    31
+1.67662657E+01+2.32109616E-02-7.93355119E-06+1.23101995E-09-7.13892514E-14    2
-2.93324539E+03-6.44104411E+01-3.63783422E-01+6.36719104E-02-4.53090160E-05    3
+1.73368393E-08-2.79133016E-12+3.04087286E+03+2.75469470E+01+0.00000000E+00    4
C6H101-5   4/12/13 THERMC   6H  10    0    0G   300.000  5000.000 1413.000    21
+1.60456030E+01+2.34774145E-02-7.85797929E-06+1.20200542E-09-6.90100029E-14    2
+2.11899382E+03-5.88452460E+01-1.01375402E+00+6.38242808E-02-4.40653860E-05    3
+1.58295163E-08-2.30830701E-12+7.94033696E+03+3.25056094E+01+0.00000000E+00    4
C6H9-A    10/17/16      C   6H   9    0    0G   300.000  5000.000 1382.000    21!CWZ NEW THERM
 1.70376899E+01 2.05549167E-02-6.96491767E-06 1.07546988E-09-6.21898909E-14    2
 1.95752798E+04-6.38078119E+01-7.24108264E-01 6.00319387E-02-3.96639738E-05    3
 1.30603563E-08-1.70075722E-12 2.59153586E+04 3.22514932E+01                   4
C6H9-A    12/ 5/12 THERMC   6H   9    0    0G   300.000  5000.000 1400.000    21
+1.70842767E+01+2.08842788E-02-7.14529004E-06+1.10943563E-09-6.43676989E-14    2
+2.01040204E+04-6.39326012E+01-2.66715213E+00+7.26196475E-02-6.05323920E-05    3
+2.66000571E-08-4.74613408E-12+2.64415017E+04+4.02220332E+01+0.00000000E+00    4
NC7H16                  C   7H  16    0    0G   300.000  5000.000 1395.000    61
+2.25012314E+01+3.46122447E-02-1.18043982E-05+1.82894500E-09-1.05955678E-13    2
-3.43062239E+04-9.33711818E+01-9.08407323E-01+8.52753530E-02-5.25668671E-05    3
+1.62954250E-08-2.01050130E-12-2.57434808E+04+3.38295611E+01+0.00000000E+00    4
C7H15-1                 C   7H  15    0    0G   300.000  5000.000 1395.000    61
+2.18654648E+01+3.27099467E-02-1.11707195E-05+1.73230780E-09-1.00418683E-13    2
-9.16995934E+03-8.64724252E+01-5.22253662E-01+8.16834621E-02-5.13242874E-05    3
+1.64263255E-08-2.12850251E-12-1.02468974E+03+3.50045259E+01+0.00000000E+00    4
C7H15-2                 C   7H  15    0    0G   300.000  5000.000 1396.000    61
+2.14174224E+01+3.28392073E-02-1.11628188E-05+1.72585155E-09-9.98390142E-14    2
-1.06455467E+04-8.35962465E+01+3.97035978E-01+7.41511374E-02-3.83235778E-05    3
+7.74076842E-09-1.21846705E-13-2.61270661E+03+3.19805516E+01+0.00000000E+00    4
C7H15-3                 C   7H  15    0    0G   300.000  5000.000 1396.000    61
+2.14174224E+01+3.28392073E-02-1.11628188E-05+1.72585155E-09-9.98390142E-14    2
-1.06455467E+04-8.35962465E+01+3.97035978E-01+7.41511374E-02-3.83235778E-05    3
+7.74076842E-09-1.21846705E-13-2.61270661E+03+3.19805516E+01+0.00000000E+00    4
C7H15-4                 C   7H  15    0    0G   300.000  5000.000 1396.000    61
+2.14174224E+01+3.28392073E-02-1.11628188E-05+1.72585155E-09-9.98390142E-14    2
-1.06455467E+04-8.42857282E+01+3.97035978E-01+7.41511374E-02-3.83235778E-05    3
+7.74076842E-09-1.21846705E-13-2.61270661E+03+3.12910700E+01+0.00000000E+00    4
C7H15OOH-1              C   7H  16O   2    0G   300.000  5000.000 1393.000    81
+2.79204752E+01+3.47496458E-02-1.19627560E-05+1.86536439E-09-1.08554328E-13    2
-4.57936217E+04-1.15336506E+02+2.44103755E-02+9.72280184E-02-6.48026839E-05    3
+2.19866894E-08-3.02783193E-12-3.58214014E+04+3.54617251E+01+0.00000000E+00    4
C7H15OOH-2              C   7H  16O   2    0G   300.000  5000.000 1400.000    81
+2.83104576E+01+3.39515981E-02-1.15841285E-05+1.79549391E-09-1.04049983E-13    2
-4.76576895E+04-1.18022294E+02+4.26850488E-01+9.92387786E-02-6.99733098E-05    3
+2.55385488E-08-3.80729481E-12-3.80148806E+04+3.16318606E+01+0.00000000E+00    4
C7H15OOH-3              C   7H  16O   2    0G   300.000  5000.000 1400.000    81
+2.83104576E+01+3.39515981E-02-1.15841285E-05+1.79549391E-09-1.04049983E-13    2
-4.76576895E+04-1.18022294E+02+4.26850488E-01+9.92387786E-02-6.99733098E-05    3
+2.55385488E-08-3.80729481E-12-3.80148806E+04+3.16318606E+01+0.00000000E+00    4
C7H15OOH-4              C   7H  16O   2    0G   300.000  5000.000 1400.000    81
+2.83104576E+01+3.39515981E-02-1.15841285E-05+1.79549391E-09-1.04049983E-13    2
-4.76576895E+04-1.18711776E+02+4.26850488E-01+9.92387786E-02-6.99733098E-05    3
+2.55385488E-08-3.80729481E-12-3.80148806E+04+3.09423790E+01+0.00000000E+00    4
C7H15-1O2               C   7H  15O   2    0G   300.000  5000.000 1392.000    71
+2.69033908E+01+3.34773175E-02-1.15204570E-05+1.79592321E-09-1.04493268E-13    2
-2.85365673E+04-1.08980069E+02+8.36337744E-01+9.12081598E-02-5.96066427E-05    3
+1.97488007E-08-2.64615990E-12-1.91440702E+04+3.21770108E+01+0.00000000E+00    4
C7H15-2O2               C   7H  15O   2    0G   300.000  5000.000 1399.000    71
+2.72644843E+01+3.26945656E-02-1.11450170E-05+1.72632915E-09-9.99959530E-14    2
-3.03857809E+04-1.11491892E+02+1.20198260E+00+9.33836346E-02-6.50845852E-05    3
+2.35152589E-08-3.47595547E-12-2.13315851E+04+2.85195439E+01+0.00000000E+00    4
C7H15-3O2               C   7H  15O   2    0G   300.000  5000.000 1399.000    71
+2.72644843E+01+3.26945656E-02-1.11450170E-05+1.72632915E-09-9.99959530E-14    2
-3.03857809E+04-1.11491892E+02+1.20198260E+00+9.33836346E-02-6.50845852E-05    3
+2.35152589E-08-3.47595547E-12-2.13315851E+04+2.85195439E+01+0.00000000E+00    4
C7H15-4O2               C   7H  15O   2    0G   300.000  5000.000 1399.000    71
+2.72644843E+01+3.26945656E-02-1.11450170E-05+1.72632915E-09-9.99959530E-14    2
-3.03857809E+04-1.12181374E+02+1.20198260E+00+9.33836346E-02-6.50845852E-05    3
+2.35152589E-08-3.47595547E-12-2.13315851E+04+2.78300623E+01+0.00000000E+00    4
C7H15-1O                C   7H  15O   1    0G   300.000  5000.000 1396.000    61
+2.54635504E+01+3.22254199E-02-1.10128382E-05+1.70895056E-09-9.91208953E-14    2
-2.68244738E+04-1.04477256E+02+1.08712676E+00+8.37177054E-02-4.99666505E-05    3
+1.38344242E-08-1.30534462E-12-1.78779963E+04+2.82643327E+01+0.00000000E+00    4
C7H15-2O                C   7H  15O   1    0G   300.000  5000.000 1404.000    61
+2.51497576E+01+3.20423962E-02-1.08501319E-05+1.67316908E-09-9.66167291E-14    2
-2.84846401E+04-1.03072531E+02+1.24372086E+00+8.52381806E-02-5.46532468E-05    3
+1.74130635E-08-2.15461900E-12-1.99857138E+04+2.61409435E+01+0.00000000E+00    4
C7H15-3O                C   7H  15O   1    0G   300.000  5000.000 1404.000    61
+2.51497576E+01+3.20423962E-02-1.08501319E-05+1.67316908E-09-9.66167291E-14    2
-2.84846401E+04-1.03072531E+02+1.24372086E+00+8.52381806E-02-5.46532468E-05    3
+1.74130635E-08-2.15461900E-12-1.99857138E+04+2.61409435E+01+0.00000000E+00    4
C7H15-4O                C   7H  15O   1    0G   300.000  5000.000 1404.000    61
+2.51497576E+01+3.20423962E-02-1.08501319E-05+1.67316908E-09-9.66167291E-14    2
-2.84846401E+04-1.03762012E+02+1.24372086E+00+8.52381806E-02-5.46532468E-05    3
+1.74130635E-08-2.15461900E-12-1.99857138E+04+2.54514619E+01+0.00000000E+00    4
C7H14OOH1-2             C   7H  15O   2    0G   300.000  5000.000 1392.000    81
+2.67171408E+01+3.31297539E-02-1.13820614E-05+1.77234804E-09-1.03039297E-13    2
-2.16844611E+04-1.05713265E+02+2.05850536E+00+8.70775096E-02-5.55512656E-05    3
+1.78824057E-08-2.31482549E-12-1.27240467E+04+2.80673449E+01+0.00000000E+00    4
C7H14OOH1-3             C   7H  15O   2    0G   300.000  5000.000 1396.000    81
+2.61247110E+01+3.33101840E-02-1.13748810E-05+1.76415357E-09-1.02280823E-13    2
-2.17289232E+04-1.01864981E+02+1.63529329E+00+8.52179548E-02-5.10436504E-05    3
+1.44161078E-08-1.44169760E-12-1.27398444E+04+3.14605052E+01+0.00000000E+00    4
C7H14OOH1-4             C   7H  15O   2    0G   300.000  5000.000 1396.000    81
+2.61247110E+01+3.33101840E-02-1.13748810E-05+1.76415357E-09-1.02280823E-13    2
-2.17289232E+04-1.01864981E+02+1.63529329E+00+8.52179548E-02-5.10436504E-05    3
+1.44161078E-08-1.44169760E-12-1.27398444E+04+3.14605052E+01+0.00000000E+00    4
C7H14OOH1-5             C   7H  15O   2    0G   300.000  5000.000 1396.000    81
+2.61247110E+01+3.33101840E-02-1.13748810E-05+1.76415357E-09-1.02280823E-13    2
-2.17289232E+04-1.01864981E+02+1.63529329E+00+8.52179548E-02-5.10436504E-05    3
+1.44161078E-08-1.44169760E-12-1.27398444E+04+3.14605052E+01+0.00000000E+00    4
C7H14OOH2-1             C   7H  15O   2    0G   300.000  5000.000 1400.000    81
+2.79788938E+01+3.17340951E-02-1.08300553E-05+1.67892063E-09-9.73081404E-14    2
-2.26191550E+04-1.13340193E+02+1.28356907E+00+9.44955667E-02-6.71910982E-05    3
+2.46830552E-08-3.69644605E-12-1.34221407E+04+2.98300713E+01+0.00000000E+00    4
C7H14OOH2-3             C   7H  15O   2    0G   300.000  5000.000 1400.000    81
+2.70174196E+01+3.23668637E-02-1.10064699E-05+1.70200278E-09-9.84688459E-14    2
-2.34973718E+04-1.07846478E+02+2.37029828E+00+8.95430479E-02-6.16372659E-05    3
+2.20878637E-08-3.24866065E-12-1.49038443E+04+2.46535755E+01+0.00000000E+00    4
C7H14OOH2-4             C   7H  15O   2    0G   300.000  5000.000 1405.000    81
+2.64783436E+01+3.24715176E-02-1.09678712E-05+1.68846547E-09-9.73849101E-14    2
-2.35623223E+04-1.04295327E+02+1.97904247E+00+8.76230614E-02-5.70967697E-05    3
+1.86207763E-08-2.37904286E-12-1.49267710E+04+2.78812322E+01+0.00000000E+00    4
C7H14OOH2-5             C   7H  15O   2    0G   300.000  5000.000 1405.000    81
+2.64783436E+01+3.24715176E-02-1.09678712E-05+1.68846547E-09-9.73849101E-14    2
-2.35623223E+04-1.04295327E+02+1.97904247E+00+8.76230614E-02-5.70967697E-05    3
+1.86207763E-08-2.37904286E-12-1.49267710E+04+2.78812322E+01+0.00000000E+00    4
C7H14OOH2-6             C   7H  15O   2    0G   300.000  5000.000 1405.000    81
+2.64783436E+01+3.24715176E-02-1.09678712E-05+1.68846547E-09-9.73849101E-14    2
-2.35623223E+04-1.04295327E+02+1.97904247E+00+8.76230614E-02-5.70967697E-05    3
+1.86207763E-08-2.37904286E-12-1.49267710E+04+2.78812322E+01+0.00000000E+00    4
C7H14OOH3-1             C   7H  15O   2    0G   300.000  5000.000 1401.000    81
+2.77319787E+01+3.19075024E-02-1.08816708E-05+1.68610984E-09-9.76912162E-14    2
-2.25232133E+04-1.12089257E+02+7.83262392E-01+9.58377482E-02-6.90031735E-05    3
+2.57734796E-08-3.93245841E-12-1.32935004E+04+3.22410995E+01+0.00000000E+00    4
C7H14OOH3-2             C   7H  15O   2    0G   300.000  5000.000 1400.000    81
+2.70174196E+01+3.23668637E-02-1.10064699E-05+1.70200278E-09-9.84688459E-14    2
-2.34973718E+04-1.07846478E+02+2.37029828E+00+8.95430479E-02-6.16372659E-05    3
+2.20878637E-08-3.24866065E-12-1.49038443E+04+2.46535755E+01+0.00000000E+00    4
C7H14OOH3-4             C   7H  15O   2    0G   300.000  5000.000 1400.000    81
+2.70174196E+01+3.23668637E-02-1.10064699E-05+1.70200278E-09-9.84688459E-14    2
-2.34973718E+04-1.07846478E+02+2.37029828E+00+8.95430479E-02-6.16372659E-05    3
+2.20878637E-08-3.24866065E-12-1.49038443E+04+2.46535755E+01+0.00000000E+00    4
C7H14OOH3-5             C   7H  15O   2    0G   300.000  5000.000 1405.000    81
+2.64783436E+01+3.24715176E-02-1.09678712E-05+1.68846547E-09-9.73849101E-14    2
-2.35623223E+04-1.04295327E+02+1.97904247E+00+8.76230614E-02-5.70967697E-05    3
+1.86207763E-08-2.37904286E-12-1.49267710E+04+2.78812322E+01+0.00000000E+00    4
C7H14OOH3-6             C   7H  15O   2    0G   300.000  5000.000 1405.000    81
+2.64783436E+01+3.24715176E-02-1.09678712E-05+1.68846547E-09-9.73849101E-14    2
-2.35623223E+04-1.04295327E+02+1.97904247E+00+8.76230614E-02-5.70967697E-05    3
+1.86207763E-08-2.37904286E-12-1.49267710E+04+2.78812322E+01+0.00000000E+00    4
C7H14OOH3-7             C   7H  15O   2    0G   300.000  5000.000 1401.000    81
+2.77319787E+01+3.19075024E-02-1.08816708E-05+1.68610984E-09-9.76912162E-14    2
-2.25232133E+04-1.12089257E+02+7.83262392E-01+9.58377482E-02-6.90031735E-05    3
+2.57734796E-08-3.93245841E-12-1.32935004E+04+3.22410995E+01+0.00000000E+00    4
C7H14OOH4-1             C   7H  15O   2    0G   300.000  5000.000 1401.000    81
+2.77319787E+01+3.19075024E-02-1.08816708E-05+1.68610984E-09-9.76912162E-14    2
-2.25232133E+04-1.12089257E+02+7.83262392E-01+9.58377482E-02-6.90031735E-05    3
+2.57734796E-08-3.93245841E-12-1.32935004E+04+3.22410995E+01+0.00000000E+00    4
C7H14OOH4-2             C   7H  15O   2    0G   300.000  5000.000 1405.000    81
+2.64783436E+01+3.24715176E-02-1.09678712E-05+1.68846547E-09-9.73849101E-14    2
-2.35623223E+04-1.04295327E+02+1.97904247E+00+8.76230614E-02-5.70967697E-05    3
+1.86207763E-08-2.37904286E-12-1.49267710E+04+2.78812322E+01+0.00000000E+00    4
C7H14OOH4-3             C   7H  15O   2    0G   300.000  5000.000 1400.000    81
+2.70174196E+01+3.23668637E-02-1.10064699E-05+1.70200278E-09-9.84688459E-14    2
-2.34973718E+04-1.07846478E+02+2.37029828E+00+8.95430479E-02-6.16372659E-05    3
+2.20878637E-08-3.24866065E-12-1.49038443E+04+2.46535755E+01+0.00000000E+00    4
C7H14O1-2               C   7H  14O   1    0G   300.000  5000.000 1414.000    51
+2.43145945E+01+3.05362342E-02-1.03132608E-05+1.58780422E-09-9.15904778E-14    2
-3.33186148E+04-1.02260982E+02-5.32362173E+00+1.03536759E-01-7.88387549E-05    3
+3.06348713E-08-4.76815463E-12-2.35540552E+04+5.53222747E+01+0.00000000E+00    4
C7H14O1-3               C   7H  14O   1    0G   300.000  5000.000 1411.000    41
+2.32391552E+01+3.18991975E-02-1.07865989E-05+1.66184086E-09-9.59019930E-14    2
-3.40230033E+04-9.80085962E+01-8.99658143E+00+1.15164182E-01-9.39167665E-05    3
+3.95269170E-08-6.68442035E-12-2.37349113E+04+7.21047219E+01+0.00000000E+00    4
C7H14O1-4               C   7H  14O   1    0G   300.000  5000.000 1411.000    31
+2.26496238E+01+3.28076656E-02-1.10970702E-05+1.71006751E-09-9.87026466E-14    2
-4.41375876E+04-9.63003234E+01-1.10425162E+01+1.19583872E-01-9.73297786E-05    3
+4.07542947E-08-6.84722710E-12-3.33740756E+04+8.15634374E+01+0.00000000E+00    4
C7H14O1-5               C   7H  14O   1    0G   300.000  5000.000 1429.000    21
+2.26509224E+01+3.23685081E-02-1.07631924E-05+1.63960080E-09-9.38766936E-14    2
-4.60716250E+04-1.00525149E+02-9.23164267E+00+1.12801180E-01-8.78296182E-05    3
+3.48128430E-08-5.48602715E-12-3.58292882E+04+6.81950662E+01+0.00000000E+00    4
C7H14O2-3               C   7H  14O   1    0G   300.000  5000.000 1420.000    51
+2.47276035E+01+2.97928117E-02-9.97261716E-06+1.52606375E-09-8.76548896E-14    2
-3.52945321E+04-1.05104871E+02-5.31868836E+00+1.06158040E-01-8.41395170E-05    3
+3.40790710E-08-5.51100667E-12-2.56598409E+04+5.37630569E+01+0.00000000E+00    4
C7H14O2-4               C   7H  14O   1    0G   300.000  5000.000 1416.000    41
+2.35365148E+01+3.12183029E-02-1.04591524E-05+1.60125267E-09-9.19956880E-14    2
-3.59381940E+04-1.00150342E+02-8.80206542E+00+1.16925403E-01-9.81273461E-05    3
+4.23712468E-08-7.30427734E-12-2.58674984E+04+6.96783672E+01+0.00000000E+00    4
C7H14O2-5               C   7H  14O   1    0G   300.000  5000.000 1417.000    31
+2.29362709E+01+3.21249586E-02-1.07666560E-05+1.64877736E-09-9.47459639E-14    2
-4.60441457E+04-9.83699162E+01-1.08488923E+01+1.21379949E-01-1.01643749E-04    3
+4.36787302E-08-7.48641956E-12-3.55071817E+04+7.91356992E+01+0.00000000E+00    4
C7H14O2-6               C   7H  14O   1    0G   300.000  5000.000 1414.000    21
+2.33853289E+01+3.24477746E-02-1.09392447E-05+1.68205180E-09-9.69385365E-14    2
-4.85465412E+04-1.06845116E+02-1.17914477E+01+1.24658462E-01-1.04127805E-04    3
+4.45024217E-08-7.58843403E-12-3.74954472E+04+7.82418086E+01+0.00000000E+00    4
C7H14O3-4               C   7H  14O   1    0G   300.000  5000.000 1420.000    51
+2.47276035E+01+2.97928117E-02-9.97261716E-06+1.52606375E-09-8.76548896E-14    2
-3.52945321E+04-1.05104871E+02-5.31868836E+00+1.06158040E-01-8.41395170E-05    3
+3.40790710E-08-5.51100667E-12-2.56598409E+04+5.37630569E+01+0.00000000E+00    4
C7H14O3-5               C   7H  14O   1    0G   300.000  5000.000 1416.000    41
+2.35365148E+01+3.12183029E-02-1.04591524E-05+1.60125267E-09-9.19956880E-14    2
-3.59381940E+04-1.00839824E+02-8.80206542E+00+1.16925403E-01-9.81273461E-05    3
+4.23712468E-08-7.30427734E-12-2.58674984E+04+6.89888856E+01+0.00000000E+00    4
C7H14OOH1-2O2           C   7H  15O   4    0G   300.000  5000.000 1394.000    91
+3.39461015E+01+3.20348143E-02-1.10936268E-05+1.73715155E-09-1.01404253E-13    2
-4.26242723E+04-1.41965954E+02+2.32043086E+00+1.02080359E-01-6.80665886E-05    3
+2.17353894E-08-2.61149960E-12-3.13880160E+04+2.90263218E+01+0.00000000E+00    4
C7H14OOH1-3O2           C   7H  15O   4    0G   300.000  5000.000 1394.000    91
+3.39461015E+01+3.20348143E-02-1.10936268E-05+1.73715155E-09-1.01404253E-13    2
-4.26242723E+04-1.41965954E+02+2.32043086E+00+1.02080359E-01-6.80665886E-05    3
+2.17353894E-08-2.61149960E-12-3.13880160E+04+2.90263218E+01+0.00000000E+00    4
C7H14OOH1-4O2           C   7H  15O   4    0G   300.000  5000.000 1394.000    91
+3.39461015E+01+3.20348143E-02-1.10936268E-05+1.73715155E-09-1.01404253E-13    2
-4.26242723E+04-1.41965954E+02+2.32043086E+00+1.02080359E-01-6.80665886E-05    3
+2.17353894E-08-2.61149960E-12-3.13880160E+04+2.90263218E+01+0.00000000E+00    4
C7H14OOH1-5O2           C   7H  15O   4    0G   300.000  5000.000 1394.000    91
+3.39461015E+01+3.20348143E-02-1.10936268E-05+1.73715155E-09-1.01404253E-13    2
-4.26242723E+04-1.41965954E+02+2.32043086E+00+1.02080359E-01-6.80665886E-05    3
+2.17353894E-08-2.61149960E-12-3.13880160E+04+2.90263218E+01+0.00000000E+00    4
C7H14OOH2-1O2           C   7H  15O   4    0G   300.000  5000.000 1394.000    91
+3.39461015E+01+3.20348143E-02-1.10936268E-05+1.73715155E-09-1.01404253E-13    2
-4.26242723E+04-1.41965954E+02+2.32043086E+00+1.02080359E-01-6.80665886E-05    3
+2.17353894E-08-2.61149960E-12-3.13880160E+04+2.90263218E+01+0.00000000E+00    4
C7H14OOH2-3O2           C   7H  15O   4    0G   300.000  5000.000 1401.000    91
+3.15622698E+01+3.32979030E-02-1.13556840E-05+1.75955945E-09-1.01947462E-13    2
-4.33174833E+04-1.28497441E+02+2.10052868E+00+1.04869368E-01-7.84344393E-05    3
+3.05606489E-08-4.86428857E-12-3.33943428E+04+2.86976000E+01+0.00000000E+00    4
C7H14OOH2-4O2           C   7H  15O   4    0G   300.000  5000.000 1401.000    91
+3.15622698E+01+3.32979030E-02-1.13556840E-05+1.75955945E-09-1.01947462E-13    2
-4.33174833E+04-1.28497441E+02+2.10052868E+00+1.04869368E-01-7.84344393E-05    3
+3.05606489E-08-4.86428857E-12-3.33943428E+04+2.86976000E+01+0.00000000E+00    4
C7H14OOH2-5O2           C   7H  15O   4    0G   300.000  5000.000 1401.000    91
+3.15622698E+01+3.32979030E-02-1.13556840E-05+1.75955945E-09-1.01947462E-13    2
-4.33174833E+04-1.28497441E+02+2.10052868E+00+1.04869368E-01-7.84344393E-05    3
+3.05606489E-08-4.86428857E-12-3.33943428E+04+2.86976000E+01+0.00000000E+00    4
C7H14OOH2-6O2           C   7H  15O   4    0G   300.000  5000.000 1401.000    91
+3.15622698E+01+3.32979030E-02-1.13556840E-05+1.75955945E-09-1.01947462E-13    2
-4.33174833E+04-1.28497441E+02+2.10052868E+00+1.04869368E-01-7.84344393E-05    3
+3.05606489E-08-4.86428857E-12-3.33943428E+04+2.86976000E+01+0.00000000E+00    4
C7H14OOH3-1O2           C   7H  15O   4    0G   300.000  5000.000 1394.000    91
+3.39461015E+01+3.20348143E-02-1.10936268E-05+1.73715155E-09-1.01404253E-13    2
-4.26242723E+04-1.41965954E+02+2.32043086E+00+1.02080359E-01-6.80665886E-05    3
+2.17353894E-08-2.61149960E-12-3.13880160E+04+2.90263218E+01+0.00000000E+00    4
C7H14OOH3-2O2           C   7H  15O   4    0G   300.000  5000.000 1401.000    91
+3.15622698E+01+3.32979030E-02-1.13556840E-05+1.75955945E-09-1.01947462E-13    2
-4.33174833E+04-1.28497441E+02+2.10052868E+00+1.04869368E-01-7.84344393E-05    3
+3.05606489E-08-4.86428857E-12-3.33943428E+04+2.86976000E+01+0.00000000E+00    4
C7H14OOH3-4O2           C   7H  15O   4    0G   300.000  5000.000 1401.000    91
+3.15622698E+01+3.32979030E-02-1.13556840E-05+1.75955945E-09-1.01947462E-13    2
-4.33174833E+04-1.28497441E+02+2.10052868E+00+1.04869368E-01-7.84344393E-05    3
+3.05606489E-08-4.86428857E-12-3.33943428E+04+2.86976000E+01+0.00000000E+00    4
C7H14OOH3-5O2           C   7H  15O   4    0G   300.000  5000.000 1401.000    91
+3.15622698E+01+3.32979030E-02-1.13556840E-05+1.75955945E-09-1.01947462E-13    2
-4.33174833E+04-1.28497441E+02+2.10052868E+00+1.04869368E-01-7.84344393E-05    3
+3.05606489E-08-4.86428857E-12-3.33943428E+04+2.86976000E+01+0.00000000E+00    4
C7H14OOH3-6O2           C   7H  15O   4    0G   300.000  5000.000 1401.000    91
+3.15622698E+01+3.32979030E-02-1.13556840E-05+1.75955945E-09-1.01947462E-13    2
-4.33174833E+04-1.28497441E+02+2.10052868E+00+1.04869368E-01-7.84344393E-05    3
+3.05606489E-08-4.86428857E-12-3.33943428E+04+2.86976000E+01+0.00000000E+00    4
C7H14OOH3-7O2           C   7H  15O   4    0G   300.000  5000.000 1394.000    91
+3.39461015E+01+3.20348143E-02-1.10936268E-05+1.73715155E-09-1.01404253E-13    2
-4.26242723E+04-1.41965954E+02+2.32043086E+00+1.02080359E-01-6.80665886E-05    3
+2.17353894E-08-2.61149960E-12-3.13880160E+04+2.90263218E+01+0.00000000E+00    4
C7H14OOH4-1O2           C   7H  15O   4    0G   300.000  5000.000 1394.000    91
+3.39461015E+01+3.20348143E-02-1.10936268E-05+1.73715155E-09-1.01404253E-13    2
-4.26242723E+04-1.41965954E+02+2.32043086E+00+1.02080359E-01-6.80665886E-05    3
+2.17353894E-08-2.61149960E-12-3.13880160E+04+2.90263218E+01+0.00000000E+00    4
C7H14OOH4-2O2           C   7H  15O   4    0G   300.000  5000.000 1401.000    91
+3.15622698E+01+3.32979030E-02-1.13556840E-05+1.75955945E-09-1.01947462E-13    2
-4.33174833E+04-1.28497441E+02+2.10052868E+00+1.04869368E-01-7.84344393E-05    3
+3.05606489E-08-4.86428857E-12-3.33943428E+04+2.86976000E+01+0.00000000E+00    4
C7H14OOH4-3O2           C   7H  15O   4    0G   300.000  5000.000 1401.000    91
+3.15622698E+01+3.32979030E-02-1.13556840E-05+1.75955945E-09-1.01947462E-13    2
-4.33174833E+04-1.28497441E+02+2.10052868E+00+1.04869368E-01-7.84344393E-05    3
+3.05606489E-08-4.86428857E-12-3.33943428E+04+2.86976000E+01+0.00000000E+00    4
C7H13Q12-3              C   7H  15O   4    0G   300.000  5000.000 1394.000    01
+3.11104496E+01+3.37811838E-02-1.16385576E-05+1.81582953E-09-1.05714699E-13    2
-3.47682853E+04-1.23525460E+02+2.55872874E+00+9.88765291E-02-6.80387144E-05    3
+2.39672496E-08-3.44171664E-12-2.46878137E+04+3.03911152E+01+0.00000000E+00    4
C7H13Q12-4              C   7H  15O   4    0G   300.000  5000.000 1407.000    01
+3.13693154E+01+3.29404356E-02-1.12115259E-05+1.73492810E-09-1.00428410E-13    2
-3.47328736E+04-1.23673782E+02+3.55376575E+00+9.74103166E-02-6.74682103E-05    3
+2.36573747E-08-3.31219515E-12-2.51150477E+04+2.57349644E+01+0.00000000E+00    4
C7H13Q12-5              C   7H  15O   4    0G   300.000  5000.000 1407.000    01
+3.13693154E+01+3.29404356E-02-1.12115259E-05+1.73492810E-09-1.00428410E-13    2
-3.47328736E+04-1.23673782E+02+3.55376575E+00+9.74103166E-02-6.74682103E-05    3
+2.36573747E-08-3.31219515E-12-2.51150477E+04+2.57349644E+01+0.00000000E+00    4
C7H13Q12-6              C   7H  15O   4    0G   300.000  5000.000 1407.000    01
+3.13693154E+01+3.29404356E-02-1.12115259E-05+1.73492810E-09-1.00428410E-13    2
-3.47328736E+04-1.23673782E+02+3.55376575E+00+9.74103166E-02-6.74682103E-05    3
+2.36573747E-08-3.31219515E-12-2.51150477E+04+2.57349644E+01+0.00000000E+00    4
C7H13Q13-2              C   7H  15O   4    0G   300.000  5000.000 1394.000    01
+3.11104496E+01+3.37811838E-02-1.16385576E-05+1.81582953E-09-1.05714699E-13    2
-3.47682853E+04-1.23525460E+02+2.55872874E+00+9.88765291E-02-6.80387144E-05    3
+2.39672496E-08-3.44171664E-12-2.46878137E+04+3.03911152E+01+0.00000000E+00    4
C7H13Q13-4              C   7H  15O   4    0G   300.000  5000.000 1394.000    01
+3.11104496E+01+3.37811838E-02-1.16385576E-05+1.81582953E-09-1.05714699E-13    2
-3.47682853E+04-1.23525460E+02+2.55872874E+00+9.88765291E-02-6.80387144E-05    3
+2.39672496E-08-3.44171664E-12-2.46878137E+04+3.03911152E+01+0.00000000E+00    4
C7H13Q13-5              C   7H  15O   4    0G   300.000  5000.000 1407.000    01
+3.13693154E+01+3.29404356E-02-1.12115259E-05+1.73492810E-09-1.00428410E-13    2
-3.47328736E+04-1.23673782E+02+3.55376575E+00+9.74103166E-02-6.74682103E-05    3
+2.36573747E-08-3.31219515E-12-2.51150477E+04+2.57349644E+01+0.00000000E+00    4
C7H13Q13-6              C   7H  15O   4    0G   300.000  5000.000 1407.000    01
+3.13693154E+01+3.29404356E-02-1.12115259E-05+1.73492810E-09-1.00428410E-13    2
-3.47328736E+04-1.23673782E+02+3.55376575E+00+9.74103166E-02-6.74682103E-05    3
+2.36573747E-08-3.31219515E-12-2.51150477E+04+2.57349644E+01+0.00000000E+00    4
C7H13Q13-7              C   7H  15O   4    0G   300.000  5000.000 1395.000    01
+3.44248733E+01+3.12441717E-02-1.08303079E-05+1.69706292E-09-9.91120837E-14    2
-3.47650019E+04-1.42631701E+02+1.89525081E+00+1.04616690E-01-7.21233992E-05    3
+2.40840687E-08-3.08867509E-12-2.33506075E+04+3.27605224E+01+0.00000000E+00    4
C7H13Q14-2              C   7H  15O   4    0G   300.000  5000.000 1394.000    01
+3.11104496E+01+3.37811838E-02-1.16385576E-05+1.81582953E-09-1.05714699E-13    2
-3.47682853E+04-1.23525460E+02+2.55872874E+00+9.88765291E-02-6.80387144E-05    3
+2.39672496E-08-3.44171664E-12-2.46878137E+04+3.03911152E+01+0.00000000E+00    4
C7H13Q14-3              C   7H  15O   4    0G   300.000  5000.000 1394.000    01
+3.11104496E+01+3.37811838E-02-1.16385576E-05+1.81582953E-09-1.05714699E-13    2
-3.47682853E+04-1.23525460E+02+2.55872874E+00+9.88765291E-02-6.80387144E-05    3
+2.39672496E-08-3.44171664E-12-2.46878137E+04+3.03911152E+01+0.00000000E+00    4
C7H13Q14-5              C   7H  15O   4    0G   300.000  5000.000 1394.000    01
+3.11104496E+01+3.37811838E-02-1.16385576E-05+1.81582953E-09-1.05714699E-13    2
-3.47682853E+04-1.23525460E+02+2.55872874E+00+9.88765291E-02-6.80387144E-05    3
+2.39672496E-08-3.44171664E-12-2.46878137E+04+3.03911152E+01+0.00000000E+00    4
C7H13Q14-6              C   7H  15O   4    0G   300.000  5000.000 1407.000    01
+3.13693154E+01+3.29404356E-02-1.12115259E-05+1.73492810E-09-1.00428410E-13    2
-3.47328736E+04-1.23673782E+02+3.55376575E+00+9.74103166E-02-6.74682103E-05    3
+2.36573747E-08-3.31219515E-12-2.51150477E+04+2.57349644E+01+0.00000000E+00    4
C7H13Q14-7              C   7H  15O   4    0G   300.000  5000.000 1395.000    01
+3.44248733E+01+3.12441717E-02-1.08303079E-05+1.69706292E-09-9.91120837E-14    2
-3.47650019E+04-1.42631701E+02+1.89525081E+00+1.04616690E-01-7.21233992E-05    3
+2.40840687E-08-3.08867509E-12-2.33506075E+04+3.27605224E+01+0.00000000E+00    4
C7H13Q15-2              C   7H  15O   4    0G   300.000  5000.000 1394.000    01
+3.11104496E+01+3.37811838E-02-1.16385576E-05+1.81582953E-09-1.05714699E-13    2
-3.47682853E+04-1.23525460E+02+2.55872874E+00+9.88765291E-02-6.80387144E-05    3
+2.39672496E-08-3.44171664E-12-2.46878137E+04+3.03911152E+01+0.00000000E+00    4
C7H13Q15-3              C   7H  15O   4    0G   300.000  5000.000 1407.000    01
+3.13693154E+01+3.29404356E-02-1.12115259E-05+1.73492810E-09-1.00428410E-13    2
-3.47328736E+04-1.23673782E+02+3.55376575E+00+9.74103166E-02-6.74682103E-05    3
+2.36573747E-08-3.31219515E-12-2.51150477E+04+2.57349644E+01+0.00000000E+00    4
C7H13Q15-4              C   7H  15O   4    0G   300.000  5000.000 1394.000    01
+3.11104496E+01+3.37811838E-02-1.16385576E-05+1.81582953E-09-1.05714699E-13    2
-3.47682853E+04-1.23525460E+02+2.55872874E+00+9.88765291E-02-6.80387144E-05    3
+2.39672496E-08-3.44171664E-12-2.46878137E+04+3.03911152E+01+0.00000000E+00    4
C7H13Q15-6              C   7H  15O   4    0G   300.000  5000.000 1394.000    01
+3.11104496E+01+3.37811838E-02-1.16385576E-05+1.81582953E-09-1.05714699E-13    2
-3.47682853E+04-1.23525460E+02+2.55872874E+00+9.88765291E-02-6.80387144E-05    3
+2.39672496E-08-3.44171664E-12-2.46878137E+04+3.03911152E+01+0.00000000E+00    4
C7H13Q15-7              C   7H  15O   4    0G   300.000  5000.000 1395.000    01
+3.44248733E+01+3.12441717E-02-1.08303079E-05+1.69706292E-09-9.91120837E-14    2
-3.47650019E+04-1.42631701E+02+1.89525081E+00+1.04616690E-01-7.21233992E-05    3
+2.40840687E-08-3.08867509E-12-2.33506075E+04+3.27605224E+01+0.00000000E+00    4
C7H13Q23-1              C   7H  15O   4    0G   300.000  5000.000 1400.000    01
+3.19365916E+01+3.26878147E-02-1.11748567E-05+1.73444372E-09-1.00611702E-13    2
-3.54856308E+04-1.28537832E+02+2.08757887E+00+1.05155888E-01-7.90124539E-05    3
+3.08131621E-08-4.89988490E-12-2.54318081E+04+3.07326377E+01+0.00000000E+00    4
C7H13Q23-4              C   7H  15O   4    0G   300.000  5000.000 1399.000    01
+3.15454850E+01+3.30379900E-02-1.12996215E-05+1.75433144E-09-1.01786375E-13    2
-3.67028604E+04-1.26588613E+02+2.95741692E+00+1.00416665E-01-7.20377682E-05    3
+2.66760295E-08-4.02711692E-12-2.68680327E+04+2.66779367E+01+0.00000000E+00    4
C7H13Q23-5              C   7H  15O   4    0G   300.000  5000.000 1416.000    01
+3.17324687E+01+3.20828367E-02-1.07959105E-05+1.65770544E-09-9.54361624E-14    2
-3.65784644E+04-1.26177142E+02+3.77629806E+00+1.00155840E-01-7.38628861E-05    3
+2.80031971E-08-4.26969253E-12-2.72782158E+04+2.27588147E+01+0.00000000E+00    4
C7H13Q23-6              C   7H  15O   4    0G   300.000  5000.000 1416.000    01
+3.17324687E+01+3.20828367E-02-1.07959105E-05+1.65770544E-09-9.54361624E-14    2
-3.65784644E+04-1.26177142E+02+3.77629806E+00+1.00155840E-01-7.38628861E-05    3
+2.80031971E-08-4.26969253E-12-2.72782158E+04+2.27588147E+01+0.00000000E+00    4
C7H13Q23-7              C   7H  15O   4    0G   300.000  5000.000 1402.000    01
+3.18911575E+01+3.26442534E-02-1.11416465E-05+1.72736491E-09-1.00122806E-13    2
-3.54199828E+04-1.28339693E+02+1.64292424E+00+1.07100207E-01-8.19867837E-05    3
+3.26301624E-08-5.28865286E-12-2.53376189E+04+3.26925968E+01+0.00000000E+00    4
C7H13Q24-1              C   7H  15O   4    0G   300.000  5000.000 1400.000    01
+3.19365916E+01+3.26878147E-02-1.11748567E-05+1.73444372E-09-1.00611702E-13    2
-3.54856308E+04-1.28537832E+02+2.08757887E+00+1.05155888E-01-7.90124539E-05    3
+3.08131621E-08-4.89988490E-12-2.54318081E+04+3.07326377E+01+0.00000000E+00    4
C7H13Q24-3              C   7H  15O   4    0G   300.000  5000.000 1399.000    01
+3.15454850E+01+3.30379900E-02-1.12996215E-05+1.75433144E-09-1.01786375E-13    2
-3.67028604E+04-1.26588613E+02+2.95741692E+00+1.00416665E-01-7.20377682E-05    3
+2.66760295E-08-4.02711692E-12-2.68680327E+04+2.66779367E+01+0.00000000E+00    4
C7H13Q24-5              C   7H  15O   4    0G   300.000  5000.000 1399.000    01
+3.15454850E+01+3.30379900E-02-1.12996215E-05+1.75433144E-09-1.01786375E-13    2
-3.67028604E+04-1.26588613E+02+2.95741692E+00+1.00416665E-01-7.20377682E-05    3
+2.66760295E-08-4.02711692E-12-2.68680327E+04+2.66779367E+01+0.00000000E+00    4
C7H13Q24-6              C   7H  15O   4    0G   300.000  5000.000 1416.000    01
+3.17324687E+01+3.20828367E-02-1.07959105E-05+1.65770544E-09-9.54361624E-14    2
-3.65784644E+04-1.26177142E+02+3.77629806E+00+1.00155840E-01-7.38628861E-05    3
+2.80031971E-08-4.26969253E-12-2.72782158E+04+2.27588147E+01+0.00000000E+00    4
C7H13Q24-7              C   7H  15O   4    0G   300.000  5000.000 1402.000    01
+3.18911575E+01+3.26442534E-02-1.11416465E-05+1.72736491E-09-1.00122806E-13    2
-3.54199828E+04-1.28339693E+02+1.64292424E+00+1.07100207E-01-8.19867837E-05    3
+3.26301624E-08-5.28865286E-12-2.53376189E+04+3.26925968E+01+0.00000000E+00    4
C7H13Q25-1              C   7H  15O   4    0G   300.000  5000.000 1400.000    01
+3.19365916E+01+3.26878147E-02-1.11748567E-05+1.73444372E-09-1.00611702E-13    2
-3.54856308E+04-1.28537832E+02+2.08757887E+00+1.05155888E-01-7.90124539E-05    3
+3.08131621E-08-4.89988490E-12-2.54318081E+04+3.07326377E+01+0.00000000E+00    4
C7H13Q25-3              C   7H  15O   4    0G   300.000  5000.000 1399.000    01
+3.15454850E+01+3.30379900E-02-1.12996215E-05+1.75433144E-09-1.01786375E-13    2
-3.67028604E+04-1.26588613E+02+2.95741692E+00+1.00416665E-01-7.20377682E-05    3
+2.66760295E-08-4.02711692E-12-2.68680327E+04+2.66779367E+01+0.00000000E+00    4
C7H13Q25-4              C   7H  15O   4    0G   300.000  5000.000 1399.000    01
+3.15454850E+01+3.30379900E-02-1.12996215E-05+1.75433144E-09-1.01786375E-13    2
-3.67028604E+04-1.26588613E+02+2.95741692E+00+1.00416665E-01-7.20377682E-05    3
+2.66760295E-08-4.02711692E-12-2.68680327E+04+2.66779367E+01+0.00000000E+00    4
C7H13Q25-6              C   7H  15O   4    0G   300.000  5000.000 1399.000    01
+3.15454850E+01+3.30379900E-02-1.12996215E-05+1.75433144E-09-1.01786375E-13    2
-3.67028604E+04-1.26588613E+02+2.95741692E+00+1.00416665E-01-7.20377682E-05    3
+2.66760295E-08-4.02711692E-12-2.68680327E+04+2.66779367E+01+0.00000000E+00    4
C7H13Q25-7              C   7H  15O   4    0G   300.000  5000.000 1402.000    01
+3.18911575E+01+3.26442534E-02-1.11416465E-05+1.72736491E-09-1.00122806E-13    2
-3.54199828E+04-1.28339693E+02+1.64292424E+00+1.07100207E-01-8.19867837E-05    3
+3.26301624E-08-5.28865286E-12-2.53376189E+04+3.26925968E+01+0.00000000E+00    4
C7H13Q26-1              C   7H  15O   4    0G   300.000  5000.000 1400.000    01
+3.19365916E+01+3.26878147E-02-1.11748567E-05+1.73444372E-09-1.00611702E-13    2
-3.54856308E+04-1.28537832E+02+2.08757887E+00+1.05155888E-01-7.90124539E-05    3
+3.08131621E-08-4.89988490E-12-2.54318081E+04+3.07326377E+01+0.00000000E+00    4
C7H13Q26-3              C   7H  15O   4    0G   300.000  5000.000 1399.000    01
+3.15454850E+01+3.30379900E-02-1.12996215E-05+1.75433144E-09-1.01786375E-13    2
-3.67028604E+04-1.26588613E+02+2.95741692E+00+1.00416665E-01-7.20377682E-05    3
+2.66760295E-08-4.02711692E-12-2.68680327E+04+2.66779367E+01+0.00000000E+00    4
C7H13Q26-4              C   7H  15O   4    0G   300.000  5000.000 1416.000    01
+3.17324687E+01+3.20828367E-02-1.07959105E-05+1.65770544E-09-9.54361624E-14    2
-3.65784644E+04-1.26866623E+02+3.77629806E+00+1.00155840E-01-7.38628861E-05    3
+2.80031971E-08-4.26969253E-12-2.72782158E+04+2.20693331E+01+0.00000000E+00    4
C7H13Q34-1              C   7H  15O   4    0G   300.000  5000.000 1402.000    01
+3.18911575E+01+3.26442534E-02-1.11416465E-05+1.72736491E-09-1.00122806E-13    2
-3.54199828E+04-1.28339693E+02+1.64292424E+00+1.07100207E-01-8.19867837E-05    3
+3.26301624E-08-5.28865286E-12-2.53376189E+04+3.26925968E+01+0.00000000E+00    4
C7H13Q34-2              C   7H  15O   4    0G   300.000  5000.000 1399.000    01
+3.15454850E+01+3.30379900E-02-1.12996215E-05+1.75433144E-09-1.01786375E-13    2
-3.67028604E+04-1.26588613E+02+2.95741692E+00+1.00416665E-01-7.20377682E-05    3
+2.66760295E-08-4.02711692E-12-2.68680327E+04+2.66779367E+01+0.00000000E+00    4
C7H13Q34-5              C   7H  15O   4    0G   300.000  5000.000 1399.000    01
+3.15454850E+01+3.30379900E-02-1.12996215E-05+1.75433144E-09-1.01786375E-13    2
-3.67028604E+04-1.26588613E+02+2.95741692E+00+1.00416665E-01-7.20377682E-05    3
+2.66760295E-08-4.02711692E-12-2.68680327E+04+2.66779367E+01+0.00000000E+00    4
C7H13Q34-6              C   7H  15O   4    0G   300.000  5000.000 1416.000    01
+3.17324687E+01+3.20828367E-02-1.07959105E-05+1.65770544E-09-9.54361624E-14    2
-3.65784644E+04-1.26177142E+02+3.77629806E+00+1.00155840E-01-7.38628861E-05    3
+2.80031971E-08-4.26969253E-12-2.72782158E+04+2.27588147E+01+0.00000000E+00    4
C7H13Q34-7              C   7H  15O   4    0G   300.000  5000.000 1402.000    01
+3.18911575E+01+3.26442534E-02-1.11416465E-05+1.72736491E-09-1.00122806E-13    2
-3.54199828E+04-1.28339693E+02+1.64292424E+00+1.07100207E-01-8.19867837E-05    3
+3.26301624E-08-5.28865286E-12-2.53376189E+04+3.26925968E+01+0.00000000E+00    4
C7H13Q35-1              C   7H  15O   4    0G   300.000  5000.000 1402.000    01
+3.18911575E+01+3.26442534E-02-1.11416465E-05+1.72736491E-09-1.00122806E-13    2
-3.54199828E+04-1.28339693E+02+1.64292424E+00+1.07100207E-01-8.19867837E-05    3
+3.26301624E-08-5.28865286E-12-2.53376189E+04+3.26925968E+01+0.00000000E+00    4
C7H13Q35-2              C   7H  15O   4    0G   300.000  5000.000 1399.000    01
+3.15454850E+01+3.30379900E-02-1.12996215E-05+1.75433144E-09-1.01786375E-13    2
-3.67028604E+04-1.26588613E+02+2.95741692E+00+1.00416665E-01-7.20377682E-05    3
+2.66760295E-08-4.02711692E-12-2.68680327E+04+2.66779367E+01+0.00000000E+00    4
C7H13Q35-4              C   7H  15O   4    0G   300.000  5000.000 1399.000    01
+3.15454850E+01+3.30379900E-02-1.12996215E-05+1.75433144E-09-1.01786375E-13    2
-3.67028604E+04-1.27278094E+02+2.95741692E+00+1.00416665E-01-7.20377682E-05    3
+2.66760295E-08-4.02711692E-12-2.68680327E+04+2.59884551E+01+0.00000000E+00    4
C7KET12                 C   7H  14O   3    0G   300.000  5000.000 1390.000    81
+3.21223692E+01+2.88333382E-02-9.97575694E-06+1.56155835E-09-9.11448835E-14    2
-5.73768969E+04-1.34951154E+02-2.02242043E+00+1.12821844E-01-8.98095474E-05    3
+3.63816839E-08-5.94859432E-12-4.60022679E+04+4.68313970E+01+0.00000000E+00    4
C7KET13                 C   7H  14O   3    0G   300.000  5000.000 1402.000    81
+2.91813264E+01+3.06159792E-02-1.04267352E-05+1.61442722E-09-9.34999392E-14    2
-5.76128277E+04-1.18979172E+02+2.41898199E+00+9.14834081E-02-6.19852852E-05    3
+2.08525236E-08-2.74537474E-12-4.82605221E+04+2.51567336E+01+0.00000000E+00    4
C7KET14                 C   7H  14O   3    0G   300.000  5000.000 1402.000    81
+2.91813264E+01+3.06159792E-02-1.04267352E-05+1.61442722E-09-9.34999392E-14    2
-5.76128277E+04-1.18979172E+02+2.41898199E+00+9.14834081E-02-6.19852852E-05    3
+2.08525236E-08-2.74537474E-12-4.82605221E+04+2.51567336E+01+0.00000000E+00    4
C7KET15                 C   7H  14O   3    0G   300.000  5000.000 1402.000    81
+2.91813264E+01+3.06159792E-02-1.04267352E-05+1.61442722E-09-9.34999392E-14    2
-5.76128277E+04-1.18979172E+02+2.41898199E+00+9.14834081E-02-6.19852852E-05    3
+2.08525236E-08-2.74537474E-12-4.82605221E+04+2.51567336E+01+0.00000000E+00    4
C7KET21                 C   7H  14O   3    0G   300.000  5000.000 1389.000    81
+3.14444661E+01+2.82938404E-02-9.56190743E-06+1.47466499E-09-8.52261942E-14    2
-5.86177087E+04-1.30228931E+02-9.11013275E-01+1.05401720E-01-7.90340286E-05    3
+2.95805586E-08-4.39236203E-12-4.77018288E+04+4.27222446E+01+0.00000000E+00    4
C7KET23                 C   7H  14O   3    0G   300.000  5000.000 1389.000    81
+3.12382757E+01+2.85248727E-02-9.65119985E-06+1.48938978E-09-8.61088842E-14    2
-6.05952490E+04-1.29479139E+02-1.30311497E+00+1.08994337E-01-8.63150634E-05    3
+3.48894872E-08-5.68162568E-12-4.98340952E+04+4.35554482E+01+0.00000000E+00    4
C7KET24                 C   7H  14O   3    0G   300.000  5000.000 1407.000    81
+2.78320035E+01+3.10208344E-02-1.04056155E-05+1.59462341E-09-9.16859524E-14    2
-6.06431441E+04-1.10882439E+02+3.08590825E+00+8.80932737E-02-5.96048275E-05    3
+2.03540139E-08-2.74781807E-12-5.20881665E+04+2.20900858E+01+0.00000000E+00    4
C7KET25                 C   7H  14O   3    0G   300.000  5000.000 1407.000    81
+2.78320035E+01+3.10208344E-02-1.04056155E-05+1.59462341E-09-9.16859524E-14    2
-6.06431441E+04-1.10882439E+02+3.08590825E+00+8.80932737E-02-5.96048275E-05    3
+2.03540139E-08-2.74781807E-12-5.20881665E+04+2.20900858E+01+0.00000000E+00    4
C7KET26                 C   7H  14O   3    0G   300.000  5000.000 1407.000    81
+2.78320035E+01+3.10208344E-02-1.04056155E-05+1.59462341E-09-9.16859524E-14    2
-6.06431441E+04-1.10882439E+02+3.08590825E+00+8.80932737E-02-5.96048275E-05    3
+2.03540139E-08-2.74781807E-12-5.20881665E+04+2.20900858E+01+0.00000000E+00    4
C7KET31                 C   7H  14O   3    0G   300.000  5000.000 1390.000    81
+2.79601586E+01+3.11058370E-02-1.04861877E-05+1.61318565E-09-9.30289704E-14    2
-5.91317971E+04-1.11897334E+02+3.35039028E+00+8.09796926E-02-4.44520581E-05    3
+9.57077658E-09-2.16392321E-13-4.99968138E+04+2.26845250E+01+0.00000000E+00    4
C7KET32                 C   7H  14O   3    0G   300.000  5000.000 1387.000    81
+3.13654946E+01+2.83825370E-02-9.59763655E-06+1.48080243E-09-8.56069968E-14    2
-6.07950743E+04-1.30969387E+02-4.64885680E-01+1.03357179E-01-7.61139823E-05    3
+2.78751565E-08-4.03730693E-12-4.99658596E+04+3.94918604E+01+0.00000000E+00    4
C7KET34                 C   7H  14O   3    0G   300.000  5000.000 1387.000    81
+3.13654946E+01+2.83825370E-02-9.59763655E-06+1.48080243E-09-8.56069968E-14    2
-6.07950743E+04-1.30969387E+02-4.64885680E-01+1.03357179E-01-7.61139823E-05    3
+2.78751565E-08-4.03730693E-12-4.99658596E+04+3.94918604E+01+0.00000000E+00    4
C7KET35                 C   7H  14O   3    0G   300.000  5000.000 1417.000    81
+2.84100629E+01+3.01275691E-02-1.00222243E-05+1.52798696E-09-8.75629841E-14    2
-6.10111353E+04-1.14884421E+02+3.76145969E+00+8.29743491E-02-4.97519839E-05    3
+1.32373155E-08-1.02452990E-12-5.21912207E+04+1.88150860E+01+0.00000000E+00    4
C7KET36                 C   7H  14O   3    0G   300.000  5000.000 1417.000    81
+2.84100629E+01+3.01275691E-02-1.00222243E-05+1.52798696E-09-8.75629841E-14    2
-6.10111353E+04-1.14884421E+02+3.76145969E+00+8.29743491E-02-4.97519839E-05    3
+1.32373155E-08-1.02452990E-12-5.21912207E+04+1.88150860E+01+0.00000000E+00    4
C7KET37                 C   7H  14O   3    0G   300.000  5000.000 1390.000    81
+2.79601586E+01+3.11058370E-02-1.04861877E-05+1.61318565E-09-9.30289704E-14    2
-5.91317971E+04-1.11897334E+02+3.35039028E+00+8.09796926E-02-4.44520581E-05    3
+9.57077658E-09-2.16392321E-13-4.99968138E+04+2.26845250E+01+0.00000000E+00    4
C7KET41                 C   7H  14O   3    0G   300.000  5000.000 1390.000    81
+2.79601586E+01+3.11058370E-02-1.04861877E-05+1.61318565E-09-9.30289704E-14    2
-5.91317971E+04-1.11897334E+02+3.35039028E+00+8.09796926E-02-4.44520581E-05    3
+9.57077658E-09-2.16392321E-13-4.99968138E+04+2.26845250E+01+0.00000000E+00    4
C7KET42                 C   7H  14O   3    0G   300.000  5000.000 1417.000    81
+2.84100629E+01+3.01275691E-02-1.00222243E-05+1.52798696E-09-8.75629841E-14    2
-6.10111353E+04-1.14884421E+02+3.76145969E+00+8.29743491E-02-4.97519839E-05    3
+1.32373155E-08-1.02452990E-12-5.21912207E+04+1.88150860E+01+0.00000000E+00    4
C7KET43                 C   7H  14O   3    0G   300.000  5000.000 1387.000    81
+3.13654946E+01+2.83825370E-02-9.59763655E-06+1.48080243E-09-8.56069968E-14    2
-6.07950743E+04-1.30969387E+02-4.64885680E-01+1.03357179E-01-7.61139823E-05    3
+2.78751565E-08-4.03730693E-12-4.99658596E+04+3.94918604E+01+0.00000000E+00    4
C7H13-1D3OOH            C   7H  14O   2    0G   300.000  5000.000 1394.000    71
+2.90779542E+01+2.88652705E-02-9.88913645E-06+1.53767589E-09-8.93288885E-14    2
-3.09726450E+04-1.22960371E+02-2.63073395E+00+1.08199467E-01-8.68167119E-05    3
+3.57892053E-08-5.96251938E-12-2.05425750E+04+4.53776182E+01+0.00000000E+00    4
C7H13-1D4OOH            C   7H  14O   2    0G   300.000  5000.000 1400.000    71
+2.62370667E+01+3.10385186E-02-1.05769230E-05+1.63789319E-09-9.48534740E-14    2
-3.13870058E+04-1.05715620E+02+7.71397342E-01+9.24620005E-02-6.79177709E-05    3
+2.62593190E-08-4.18178337E-12-2.27326381E+04+3.03693290E+01+0.00000000E+00    4
C7H13-1D5OOH            C   7H  14O   2    0G   300.000  5000.000 1400.000    71
+2.62370667E+01+3.10385186E-02-1.05769230E-05+1.63789319E-09-9.48534740E-14    2
-3.13870058E+04-1.05715620E+02+7.71397342E-01+9.24620005E-02-6.79177709E-05    3
+2.62593190E-08-4.18178337E-12-2.27326381E+04+3.03693290E+01+0.00000000E+00    4
C7H13-1D6OOH            C   7H  14O   2    0G   300.000  5000.000 1400.000    71
+2.62370667E+01+3.10385186E-02-1.05769230E-05+1.63789319E-09-9.48534740E-14    2
-3.13870058E+04-1.05715620E+02+7.71397342E-01+9.24620005E-02-6.79177709E-05    3
+2.62593190E-08-4.18178337E-12-2.27326381E+04+3.03693290E+01+0.00000000E+00    4
C7H13-2D1OOH            C   7H  14O   2    0G   300.000  5000.000 1387.000    71
+2.76028881E+01+3.04944644E-02-1.05308927E-05+1.64588437E-09-9.59461833E-14    2
-2.98877195E+04-1.12572059E+02-1.03739963E-01+9.52952380E-02-6.91621723E-05    3
+2.61655996E-08-4.09598961E-12-2.02211307E+04+3.62929671E+01+0.00000000E+00    4
C7H13-2D4OOH            C   7H  14O   2    0G   300.000  5000.000 1392.000    71
+2.87054975E+01+2.90956441E-02-9.95173224E-06+1.54585405E-09-8.97456708E-14    2
-3.21955351E+04-1.21533069E+02-1.86598369E+00+1.03608595E-01-7.99220598E-05    3
+3.16229589E-08-5.06942228E-12-2.19482737E+04+4.14584607E+01+0.00000000E+00    4
C7H13-2D5OOH            C   7H  14O   2    0G   300.000  5000.000 1399.000    71
+2.57999207E+01+3.13359785E-02-1.06638378E-05+1.64987512E-09-9.54885493E-14    2
-3.25697474E+04-1.03891031E+02+1.56048081E+00+8.78913800E-02-6.11946460E-05    3
+2.22475016E-08-3.32765732E-12-2.41452632E+04+2.63118291E+01+0.00000000E+00    4
C7H13-2D6OOH            C   7H  14O   2    0G   300.000  5000.000 1399.000    71
+2.57999207E+01+3.13359785E-02-1.06638378E-05+1.64987512E-09-9.54885493E-14    2
-3.25697474E+04-1.03891031E+02+1.56048081E+00+8.78913800E-02-6.11946460E-05    3
+2.22475016E-08-3.32765732E-12-2.41452632E+04+2.63118291E+01+0.00000000E+00    4
C7H13-2D7OOH            C   7H  14O   2    0G   300.000  5000.000 1391.000    71
+2.54707867E+01+3.21318886E-02-1.10527598E-05+1.72250760E-09-1.00200663E-13    2
-3.07525576E+04-1.01606636E+02+1.21017968E+00+8.55196199E-02-5.52653305E-05    3
+1.81653282E-08-2.42677675E-12-2.19569963E+04+2.99229828E+01+0.00000000E+00    4
C7H13-3D1OOH            C   7H  14O   2    0G   300.000  5000.000 1390.000    71
+2.51298151E+01+3.24123329E-02-1.11475843E-05+1.73711843E-09-1.01043971E-13    2
-3.06454833E+04-9.98270039E+01+8.82027682E-01+8.55388349E-02-5.48810116E-05    3
+1.78755251E-08-2.36265653E-12-2.18276358E+04+3.17219563E+01+0.00000000E+00    4
C7H13-3D2OOH            C   7H  14O   2    0G   300.000  5000.000 1390.000    71
+2.85979916E+01+2.90024472E-02-9.88429804E-06+1.53207421E-09-8.88244781E-14    2
-3.21807608E+04-1.21066515E+02-2.23029288E+00+1.03631041E-01-7.92640337E-05    3
+3.09828829E-08-4.89738221E-12-2.18100535E+04+4.34531959E+01+0.00000000E+00    4
C7H13-3D5OOH            C   7H  14O   2    0G   300.000  5000.000 1390.000    71
+2.85979916E+01+2.90024472E-02-9.88429804E-06+1.53207421E-09-8.88244781E-14    2
-3.21807608E+04-1.21066515E+02-2.23029288E+00+1.03631041E-01-7.92640337E-05    3
+3.09828829E-08-4.89738221E-12-2.18100535E+04+4.34531959E+01+0.00000000E+00    4
C7H13-3D6OOH            C   7H  14O   2    0G   300.000  5000.000 1398.000    71
+2.54729557E+01+3.16019436E-02-1.07532892E-05+1.66362284E-09-9.62810785E-14    2
-3.24718124E+04-1.02199028E+02+1.18744278E+00+8.80721168E-02-6.10131641E-05    3
+2.20696430E-08-3.28659463E-12-2.40081173E+04+2.83264595E+01+0.00000000E+00    4
C7H13-3D7OOH            C   7H  14O   2    0G   300.000  5000.000 1390.000    71
+2.51298151E+01+3.24123329E-02-1.11475843E-05+1.73711843E-09-1.01043971E-13    2
-3.06454833E+04-9.98270039E+01+8.82027682E-01+8.55388349E-02-5.48810116E-05    3
+1.78755251E-08-2.36265653E-12-2.18276358E+04+3.17219563E+01+0.00000000E+00    4
C7H13O12-3OOH           C   7H  14O   3    0G   300.000  5000.000 1423.000    71
+3.06568109E+01+2.92778514E-02-9.86078739E-06+1.51586516E-09-8.73673279E-14    2
-4.68701203E+04-1.30596042E+02-2.32721619E+00+1.10522706E-01-8.53554175E-05    3
+3.28439542E-08-4.97162723E-12-3.60936612E+04+4.46258578E+01+0.00000000E+00    4
C7H13O12-4OOH           C   7H  14O   3    0G   300.000  5000.000 1423.000    71
+3.06568109E+01+2.92778514E-02-9.86078739E-06+1.51586516E-09-8.73673279E-14    2
-4.68701203E+04-1.30596042E+02-2.32721619E+00+1.10522706E-01-8.53554175E-05    3
+3.28439542E-08-4.97162723E-12-3.60936612E+04+4.46258578E+01+0.00000000E+00    4
C7H13O12-5OOH           C   7H  14O   3    0G   300.000  5000.000 1423.000    71
+3.06568109E+01+2.92778514E-02-9.86078739E-06+1.51586516E-09-8.73673279E-14    2
-4.68701203E+04-1.30596042E+02-2.32721619E+00+1.10522706E-01-8.53554175E-05    3
+3.28439542E-08-4.97162723E-12-3.60936612E+04+4.46258578E+01+0.00000000E+00    4
C7H13O12-6OOH           C   7H  14O   3    0G   300.000  5000.000 1423.000    71
+3.06568109E+01+2.92778514E-02-9.86078739E-06+1.51586516E-09-8.73673279E-14    2
-4.68701203E+04-1.30596042E+02-2.32721619E+00+1.10522706E-01-8.53554175E-05    3
+3.28439542E-08-4.97162723E-12-3.60936612E+04+4.46258578E+01+0.00000000E+00    4
C7H13O13-2OOH           C   7H  14O   3    0G   300.000  5000.000 1420.000    61
+2.95844365E+01+3.05756089E-02-1.02984950E-05+1.58302884E-09-9.12273949E-14    2
-4.75700916E+04-1.26331319E+02-5.09972940E+00+1.17940417E-01-9.39654580E-05    3
+3.76366993E-08-5.96942332E-12-3.64053536E+04+5.72799707E+01+0.00000000E+00    4
C7H13O13-4OOH           C   7H  14O   3    0G   300.000  5000.000 1420.000    61
+2.95844365E+01+3.05756089E-02-1.02984950E-05+1.58302884E-09-9.12273949E-14    2
-4.75700916E+04-1.26331319E+02-5.09972940E+00+1.17940417E-01-9.39654580E-05    3
+3.76366993E-08-5.96942332E-12-3.64053536E+04+5.72799707E+01+0.00000000E+00    4
C7H13O13-5OOH           C   7H  14O   3    0G   300.000  5000.000 1420.000    61
+2.95844365E+01+3.05756089E-02-1.02984950E-05+1.58302884E-09-9.12273949E-14    2
-4.75700916E+04-1.26331319E+02-5.09972940E+00+1.17940417E-01-9.39654580E-05    3
+3.76366993E-08-5.96942332E-12-3.64053536E+04+5.72799707E+01+0.00000000E+00    4
C7H13O13-6OOH           C   7H  14O   3    0G   300.000  5000.000 1420.000    61
+2.95844365E+01+3.05756089E-02-1.02984950E-05+1.58302884E-09-9.12273949E-14    2
-4.75700916E+04-1.26331319E+02-5.09972940E+00+1.17940417E-01-9.39654580E-05    3
+3.76366993E-08-5.96942332E-12-3.64053536E+04+5.72799707E+01+0.00000000E+00    4
C7H13O13-7OOH           C   7H  14O   3    0G   300.000  5000.000 1426.000    61
+2.97373561E+01+3.06836196E-02-1.03914057E-05+1.60356739E-09-9.26750590E-14    2
-4.59445681E+04-1.26820023E+02-6.07792808E+00+1.17208958E-01-8.86164334E-05    3
+3.28978179E-08-4.74711308E-12-3.40965125E+04+6.40055015E+01+0.00000000E+00    4
C7H13O14-2OOH           C   7H  14O   3    0G   300.000  5000.000 1420.000    51
+2.89220143E+01+3.15527403E-02-1.06334605E-05+1.63510994E-09-9.42520946E-14    2
-5.76473124E+04-1.24190446E+02-7.38516052E+00+1.23530656E-01-9.93379244E-05    3
+4.01682077E-08-6.43221166E-12-4.60102633E+04+6.78304029E+01+0.00000000E+00    4
C7H13O14-3OOH           C   7H  14O   3    0G   300.000  5000.000 1420.000    51
+2.89220143E+01+3.15527403E-02-1.06334605E-05+1.63510994E-09-9.42520946E-14    2
-5.76473124E+04-1.24190446E+02-7.38516052E+00+1.23530656E-01-9.93379244E-05    3
+4.01682077E-08-6.43221166E-12-4.60102633E+04+6.78304029E+01+0.00000000E+00    4
C7H13O14-5OOH           C   7H  14O   3    0G   300.000  5000.000 1420.000    51
+2.89220143E+01+3.15527403E-02-1.06334605E-05+1.63510994E-09-9.42520946E-14    2
-5.76473124E+04-1.24190446E+02-7.38516052E+00+1.23530656E-01-9.93379244E-05    3
+4.01682077E-08-6.43221166E-12-4.60102633E+04+6.78304029E+01+0.00000000E+00    4
C7H13O14-6OOH           C   7H  14O   3    0G   300.000  5000.000 1420.000    51
+2.89220143E+01+3.15527403E-02-1.06334605E-05+1.63510994E-09-9.42520946E-14    2
-5.76473124E+04-1.24190446E+02-7.38516052E+00+1.23530656E-01-9.93379244E-05    3
+4.01682077E-08-6.43221166E-12-4.60102633E+04+6.78304029E+01+0.00000000E+00    4
C7H13O14-7OOH           C   7H  14O   3    0G   300.000  5000.000 1411.000    51
+2.78208253E+01+3.28577038E-02-1.11593341E-05+1.72461553E-09-9.97496498E-14    2
-5.53881549E+04-1.17204730E+02-9.47844518E+00+1.29744960E-01-1.08213683E-04    3
+4.59800558E-08-7.79516037E-12-4.35716314E+04+7.93825063E+01+0.00000000E+00    4
C7H13O15-2OOH           C   7H  14O   3    0G   300.000  5000.000 1413.000    41
+2.89783260E+01+3.22434242E-02-1.09366600E-05+1.68885807E-09-9.76309782E-14    2
-5.99348988E+04-1.29616717E+02-9.62798776E+00+1.33413575E-01-1.13026808E-04    3
+4.84924849E-08-8.26487244E-12-4.78194095E+04+7.35004874E+01+0.00000000E+00    4
C7H13O15-3OOH           C   7H  14O   3    0G   300.000  5000.000 1413.000    41
+2.89783260E+01+3.22434242E-02-1.09366600E-05+1.68885807E-09-9.76309782E-14    2
-5.99348988E+04-1.29616717E+02-9.62798776E+00+1.33413575E-01-1.13026808E-04    3
+4.84924849E-08-8.26487244E-12-4.78194095E+04+7.35004874E+01+0.00000000E+00    4
C7H13O15-4OOH           C   7H  14O   3    0G   300.000  5000.000 1413.000    41
+2.89783260E+01+3.22434242E-02-1.09366600E-05+1.68885807E-09-9.76309782E-14    2
-5.99348988E+04-1.29616717E+02-9.62798776E+00+1.33413575E-01-1.13026808E-04    3
+4.84924849E-08-8.26487244E-12-4.78194095E+04+7.35004874E+01+0.00000000E+00    4
C7H13O15-6OOH           C   7H  14O   3    0G   300.000  5000.000 1413.000    41
+2.89783260E+01+3.22434242E-02-1.09366600E-05+1.68885807E-09-9.76309782E-14    2
-5.99348988E+04-1.29616717E+02-9.62798776E+00+1.33413575E-01-1.13026808E-04    3
+4.84924849E-08-8.26487244E-12-4.78194095E+04+7.35004874E+01+0.00000000E+00    4
C7H13O15-7OOH           C   7H  14O   3    0G   300.000  5000.000 1424.000    41
+2.77068460E+01+3.25453847E-02-1.08747736E-05+1.66236264E-09-9.54208828E-14    2
-5.73018452E+04-1.20830748E+02-8.20175654E+00+1.24849412E-01-1.01351038E-04    3
+4.16384416E-08-6.78332664E-12-4.59311487E+04+6.85988386E+01+0.00000000E+00    4
C7H13O23-1OOH           C   7H  14O   3    0G   300.000  5000.000 1418.000    71
+3.00568523E+01+2.97967943E-02-1.00386897E-05+1.54327355E-09-8.89410623E-14    2
-4.66455239E+04-1.26998202E+02-3.48236315E+00+1.14929716E-01-9.24757732E-05    3
+3.75714951E-08-6.06093263E-12-3.58960850E+04+5.03515097E+01+0.00000000E+00    4
C7H13O23-4OOH           C   7H  14O   3    0G   300.000  5000.000 1430.000    71
+3.12297761E+01+2.84059813E-02-9.47956084E-06+1.44833421E-09-8.31213006E-14    2
-4.89319218E+04-1.34405365E+02-2.38926773E+00+1.13321280E-01-9.05926994E-05    3
+3.61165874E-08-5.65964024E-12-3.81876031E+04+4.33940193E+01+0.00000000E+00    4
C7H13O23-5OOH           C   7H  14O   3    0G   300.000  5000.000 1430.000    71
+3.12297761E+01+2.84059813E-02-9.47956084E-06+1.44833421E-09-8.31213006E-14    2
-4.89319218E+04-1.34405365E+02-2.38926773E+00+1.13321280E-01-9.05926994E-05    3
+3.61165874E-08-5.65964024E-12-3.81876031E+04+4.33940193E+01+0.00000000E+00    4
C7H13O23-6OOH           C   7H  14O   3    0G   300.000  5000.000 1430.000    71
+3.12297761E+01+2.84059813E-02-9.47956084E-06+1.44833421E-09-8.31213006E-14    2
-4.89319218E+04-1.34405365E+02-2.38926773E+00+1.13321280E-01-9.05926994E-05    3
+3.61165874E-08-5.65964024E-12-3.81876031E+04+4.33940193E+01+0.00000000E+00    4
C7H13O23-7OOH           C   7H  14O   3    0G   300.000  5000.000 1418.000    71
+3.00568523E+01+2.97967943E-02-1.00386897E-05+1.54327355E-09-8.89410623E-14    2
-4.66455239E+04-1.26998202E+02-3.48236315E+00+1.14929716E-01-9.24757732E-05    3
+3.75714951E-08-6.06093263E-12-3.58960850E+04+5.03515097E+01+0.00000000E+00    4
C7H13O24-1OOH           C   7H  14O   3    0G   300.000  5000.000 1418.000    61
+2.91867544E+01+3.09303975E-02-1.04230990E-05+1.60259046E-09-9.23672529E-14    2
-4.74452970E+04-1.23929207E+02-5.67998134E+00+1.19707498E-01-9.67220537E-05    3
+3.94860496E-08-6.40186846E-12-3.62950216E+04+6.03473723E+01+0.00000000E+00    4
C7H13O24-3OOH           C   7H  14O   3    0G   300.000  5000.000 1426.000    61
+3.00847400E+01+2.97514366E-02-9.93001694E-06+1.51705678E-09-8.70533351E-14    2
-4.95919063E+04-1.29697889E+02-5.12505465E+00+1.20631654E-01-9.92122912E-05    3
+4.09823768E-08-6.68221982E-12-3.85055230E+04+5.58707111E+01+0.00000000E+00    4
C7H13O24-5OOH           C   7H  14O   3    0G   300.000  5000.000 1426.000    61
+3.00847400E+01+2.97514366E-02-9.93001694E-06+1.51705678E-09-8.70533351E-14    2
-4.95919063E+04-1.29697889E+02-5.12505465E+00+1.20631654E-01-9.92122912E-05    3
+4.09823768E-08-6.68221982E-12-3.85055230E+04+5.58707111E+01+0.00000000E+00    4
C7H13O24-6OOH           C   7H  14O   3    0G   300.000  5000.000 1426.000    61
+3.00847400E+01+2.97514366E-02-9.93001694E-06+1.51705678E-09-8.70533351E-14    2
-4.95919063E+04-1.29697889E+02-5.12505465E+00+1.20631654E-01-9.92122912E-05    3
+4.09823768E-08-6.68221982E-12-3.85055230E+04+5.58707111E+01+0.00000000E+00    4
C7H13O24-7OOH           C   7H  14O   3    0G   300.000  5000.000 1418.000    61
+2.91867544E+01+3.09303975E-02-1.04230990E-05+1.60259046E-09-9.23672529E-14    2
-4.74452970E+04-1.23929207E+02-5.67998134E+00+1.19707498E-01-9.67220537E-05    3
+3.94860496E-08-6.40186846E-12-3.62950216E+04+6.03473723E+01+0.00000000E+00    4
C7H13O25-1OOH           C   7H  14O   3    0G   300.000  5000.000 1415.000    51
+2.81263101E+01+3.21834697E-02-1.08370884E-05+1.66513411E-09-9.59194966E-14    2
-5.73112488E+04-1.19400460E+02-9.35219725E+00+1.31786584E-01-1.12805010E-04    3
+4.90506384E-08-8.46416378E-12-4.56933874E+04+7.72815674E+01+0.00000000E+00    4
C7H13O25-3OOH           C   7H  14O   3    0G   300.000  5000.000 1426.000    51
+2.93895989E+01+3.07437385E-02-1.02672480E-05+1.56916906E-09-9.00663946E-14    2
-5.96489796E+04-1.27352802E+02-7.41940814E+00+1.26301646E-01-1.04795872E-04    3
+4.36768367E-08-7.18457779E-12-4.81097554E+04+6.64562231E+01+0.00000000E+00    4
C7H13O25-4OOH           C   7H  14O   3    0G   300.000  5000.000 1426.000    51
+2.93895989E+01+3.07437385E-02-1.02672480E-05+1.56916906E-09-9.00663946E-14    2
-5.96489796E+04-1.27352802E+02-7.41940814E+00+1.26301646E-01-1.04795872E-04    3
+4.36768367E-08-7.18457779E-12-4.81097554E+04+6.64562231E+01+0.00000000E+00    4
C7H13O25-6OOH           C   7H  14O   3    0G   300.000  5000.000 1426.000    51
+2.93895989E+01+3.07437385E-02-1.02672480E-05+1.56916906E-09-9.00663946E-14    2
-5.96489796E+04-1.27352802E+02-7.41940814E+00+1.26301646E-01-1.04795872E-04    3
+4.36768367E-08-7.18457779E-12-4.81097554E+04+6.64562231E+01+0.00000000E+00    4
C7H13O25-7OOH           C   7H  14O   3    0G   300.000  5000.000 1415.000    51
+2.81263101E+01+3.21834697E-02-1.08370884E-05+1.66513411E-09-9.59194966E-14    2
-5.73112488E+04-1.19400460E+02-9.35219725E+00+1.31786584E-01-1.12805010E-04    3
+4.90506384E-08-8.46416378E-12-4.56933874E+04+7.72815674E+01+0.00000000E+00    4
C7H13O26-1OOH           C   7H  14O   3    0G   300.000  5000.000 1413.000    41
+2.86273198E+01+3.24610451E-02-1.09938875E-05+1.69592937E-09-9.79672635E-14    2
-5.98085835E+04-1.27424180E+02-9.81319024E+00+1.33459969E-01-1.13207306E-04    3
+4.86930651E-08-8.32140331E-12-4.77700612E+04+7.47294038E+01+0.00000000E+00    4
C7H13O26-3OOH           C   7H  14O   3    0G   300.000  5000.000 1417.000    41
+2.93182689E+01+3.15493166E-02-1.06099989E-05+1.62896879E-09-9.37892837E-14    2
-6.18764814E+04-1.32025719E+02-9.49984301E+00+1.35464135E-01-1.17595961E-04    3
+5.15396865E-08-8.92847088E-12-4.99422805E+04+7.13802548E+01+0.00000000E+00    4
C7H13O26-4OOH           C   7H  14O   3    0G   300.000  5000.000 1417.000    41
+2.93182689E+01+3.15493166E-02-1.06099989E-05+1.62896879E-09-9.37892837E-14    2
-6.18764814E+04-1.32715201E+02-9.49984301E+00+1.35464135E-01-1.17595961E-04    3
+5.15396865E-08-8.92847088E-12-4.99422805E+04+7.06907732E+01+0.00000000E+00    4
C7H13O34-1OOH           C   7H  14O   3    0G   300.000  5000.000 1418.000    71
+3.00568523E+01+2.97967943E-02-1.00386897E-05+1.54327355E-09-8.89410623E-14    2
-4.66455239E+04-1.26998202E+02-3.48236315E+00+1.14929716E-01-9.24757732E-05    3
+3.75714951E-08-6.06093263E-12-3.58960850E+04+5.03515097E+01+0.00000000E+00    4
C7H13O34-2OOH           C   7H  14O   3    0G   300.000  5000.000 1430.000    71
+3.12297761E+01+2.84059813E-02-9.47956084E-06+1.44833421E-09-8.31213006E-14    2
-4.89319218E+04-1.34405365E+02-2.38926773E+00+1.13321280E-01-9.05926994E-05    3
+3.61165874E-08-5.65964024E-12-3.81876031E+04+4.33940193E+01+0.00000000E+00    4
C7H13O34-5OOH           C   7H  14O   3    0G   300.000  5000.000 1430.000    71
+3.12297761E+01+2.84059813E-02-9.47956084E-06+1.44833421E-09-8.31213006E-14    2
-4.89319218E+04-1.34405365E+02-2.38926773E+00+1.13321280E-01-9.05926994E-05    3
+3.61165874E-08-5.65964024E-12-3.81876031E+04+4.33940193E+01+0.00000000E+00    4
C7H13O34-6OOH           C   7H  14O   3    0G   300.000  5000.000 1430.000    71
+3.12297761E+01+2.84059813E-02-9.47956084E-06+1.44833421E-09-8.31213006E-14    2
-4.89319218E+04-1.34405365E+02-2.38926773E+00+1.13321280E-01-9.05926994E-05    3
+3.61165874E-08-5.65964024E-12-3.81876031E+04+4.33940193E+01+0.00000000E+00    4
C7H13O34-7OOH           C   7H  14O   3    0G   300.000  5000.000 1418.000    71
+3.00568523E+01+2.97967943E-02-1.00386897E-05+1.54327355E-09-8.89410623E-14    2
-4.66455239E+04-1.26998202E+02-3.48236315E+00+1.14929716E-01-9.24757732E-05    3
+3.75714951E-08-6.06093263E-12-3.58960850E+04+5.03515097E+01+0.00000000E+00    4
C7H13O35-1OOH           C   7H  14O   3    0G   300.000  5000.000 1418.000    61
+2.91867544E+01+3.09303975E-02-1.04230990E-05+1.60259046E-09-9.23672529E-14    2
-4.74452970E+04-1.23929207E+02-5.67998134E+00+1.19707498E-01-9.67220537E-05    3
+3.94860496E-08-6.40186846E-12-3.62950216E+04+6.03473723E+01+0.00000000E+00    4
C7H13O35-2OOH           C   7H  14O   3    0G   300.000  5000.000 1426.000    61
+3.00847400E+01+2.97514366E-02-9.93001694E-06+1.51705678E-09-8.70533351E-14    2
-4.95919063E+04-1.29697889E+02-5.12505465E+00+1.20631654E-01-9.92122912E-05    3
+4.09823768E-08-6.68221982E-12-3.85055230E+04+5.58707111E+01+0.00000000E+00    4
C7H13O35-4OOH           C   7H  14O   3    0G   300.000  5000.000 1426.000    61
+3.00847400E+01+2.97514366E-02-9.93001694E-06+1.51705678E-09-8.70533351E-14    2
-4.95919063E+04-1.30387371E+02-5.12505465E+00+1.20631654E-01-9.92122912E-05    3
+4.09823768E-08-6.68221982E-12-3.85055230E+04+5.51812295E+01+0.00000000E+00    4
C7KET12O                C   7H  13O   2    0G   300.000  5000.000 1383.000    61
+2.78249579E+01+2.86775775E-02-1.00138821E-05+1.57662822E-09-9.23773712E-14    2
-3.89317108E+04-1.14577628E+02+2.14339924E+00+8.14112315E-02-4.80755304E-05    3
+1.24299598E-08-9.55786972E-13-2.93375207E+04+2.58408223E+01+0.00000000E+00    4
C7KET13O                C   7H  13O   2    0G   300.000  5000.000 1393.000    61
+2.60215737E+01+2.93374256E-02-1.00488420E-05+1.56203531E-09-9.07167677E-14    2
-3.87867271E+04-1.04825481E+02+2.80462854E+00+7.58170916E-02-4.12532654E-05    3
+8.70139631E-09-1.64177572E-13-3.00690471E+04+2.24125766E+01+0.00000000E+00    4
C7KET14O                C   7H  13O   2    0G   300.000  5000.000 1393.000    61
+2.60215737E+01+2.93374256E-02-1.00488420E-05+1.56203531E-09-9.07167677E-14    2
-3.87867271E+04-1.04825481E+02+2.80462854E+00+7.58170916E-02-4.12532654E-05    3
+8.70139631E-09-1.64177572E-13-3.00690471E+04+2.24125766E+01+0.00000000E+00    4
C7KET15O                C   7H  13O   2    0G   300.000  5000.000 1393.000    61
+2.60215737E+01+2.93374256E-02-1.00488420E-05+1.56203531E-09-9.07167677E-14    2
-3.87867271E+04-1.04825481E+02+2.80462854E+00+7.58170916E-02-4.12532654E-05    3
+8.70139631E-09-1.64177572E-13-3.00690471E+04+2.24125766E+01+0.00000000E+00    4
C7KET21O                C   7H  13O   2    0G   300.000  5000.000 1554.000    61
+2.54344050E+01+2.95193155E-02-1.00512410E-05+1.55686735E-09-9.02141987E-14    2
-3.93052035E+04-1.00417355E+02+7.08469593E+00+5.76449309E-02-1.67872461E-05    3
-5.15289018E-09+2.66912467E-12-3.15428673E+04+3.22374729E+00+0.00000000E+00    4
C7KET23O                C   7H  13O   2    0G   300.000  5000.000 1389.000    61
+2.54534371E+01+3.00869490E-02-1.03619417E-05+1.61623343E-09-9.40768952E-14    2
-4.15102413E+04-1.00518430E+02+3.16633176E+00+7.66586596E-02-4.55096741E-05    3
+1.27504840E-08-1.28364522E-12-3.32138551E+04+2.11371718E+01+0.00000000E+00    4
C7KET24O                C   7H  13O   2    0G   300.000  5000.000 1424.000    61
+2.52611368E+01+2.89653302E-02-9.70051521E-06+1.48514450E-09-8.53401253E-14    2
-4.18462987E+04-9.96610355E+01+4.04551808E+00+7.28475517E-02-4.06939129E-05    3
+9.42771341E-09-4.15988455E-13-3.40727262E+04+1.60209312E+01+0.00000000E+00    4
C7KET25O                C   7H  13O   2    0G   300.000  5000.000 1424.000    61
+2.52611368E+01+2.89653302E-02-9.70051521E-06+1.48514450E-09-8.53401253E-14    2
-4.18462987E+04-9.96610355E+01+4.04551808E+00+7.28475517E-02-4.06939129E-05    3
+9.42771341E-09-4.15988455E-13-3.40727262E+04+1.60209312E+01+0.00000000E+00    4
C7KET26O                C   7H  13O   2    0G   300.000  5000.000 1424.000    61
+2.52611368E+01+2.89653302E-02-9.70051521E-06+1.48514450E-09-8.53401253E-14    2
-4.18462987E+04-9.96610355E+01+4.04551808E+00+7.28475517E-02-4.06939129E-05    3
+9.42771341E-09-4.15988455E-13-3.40727262E+04+1.60209312E+01+0.00000000E+00    4
C7KET31O                C   7H  13O   2    0G   300.000  5000.000 1404.000    61
+2.54336685E+01+2.89559213E-02-9.73523973E-06+1.49510786E-09-8.61222040E-14    2
-4.02596015E+04-1.00920853E+02+4.86648027E+00+6.45174583E-02-2.45246679E-05    3
-1.77081536E-09+2.18648284E-12-3.20963786E+04+1.35846460E+01+0.00000000E+00    4
C7KET32O                C   7H  13O   2    0G   300.000  5000.000 1387.000    61
+2.52474702E+01+3.00387223E-02-1.02980700E-05+1.60151220E-09-9.30327317E-14    2
-4.15079135E+04-9.99196024E+01+4.22370120E+00+7.02977244E-02-3.51511137E-05    3
+5.96766285E-09+2.70620719E-13-3.33805928E+04+1.60319393E+01+0.00000000E+00    4
C7KET34O                C   7H  13O   2    0G   300.000  5000.000 1387.000    61
+2.52474702E+01+3.00387223E-02-1.02980700E-05+1.60151220E-09-9.30327317E-14    2
-4.15079135E+04-9.99196024E+01+4.22370120E+00+7.02977244E-02-3.51511137E-05    3
+5.96766285E-09+2.70620719E-13-3.33805928E+04+1.60319393E+01+0.00000000E+00    4
C7KET35O                C   7H  13O   2    0G   300.000  5000.000 1370.000    61
+2.56884614E+01+2.80095890E-02-9.25680532E-06+1.40530115E-09-8.03019698E-14    2
-4.20976441E+04-1.01960623E+02+4.70018599E+00+6.81280965E-02-3.21429326E-05    3
+3.33860657E-09+1.05751924E-12-3.41777201E+04+1.34845759E+01+0.00000000E+00    4
C7KET36O                C   7H  13O   2    0G   300.000  5000.000 1370.000    61
+2.56884614E+01+2.80095890E-02-9.25680532E-06+1.40530115E-09-8.03019698E-14    2
-4.20976441E+04-1.02650105E+02+4.70018599E+00+6.81280965E-02-3.21429326E-05    3
+3.33860657E-09+1.05751924E-12-3.41777201E+04+1.27950943E+01+0.00000000E+00    4
C7KET37O                C   7H  13O   2    0G   300.000  5000.000 1404.000    61
+2.54336685E+01+2.89559213E-02-9.73523973E-06+1.49510786E-09-8.61222040E-14    2
-4.02596015E+04-1.00920853E+02+4.86648027E+00+6.45174583E-02-2.45246679E-05    3
-1.77081536E-09+2.18648284E-12-3.20963786E+04+1.35846460E+01+0.00000000E+00    4
C7KET41O                C   7H  13O   2    0G   300.000  5000.000 1404.000    61
+2.54336685E+01+2.89559213E-02-9.73523973E-06+1.49510786E-09-8.61222040E-14    2
-4.02596015E+04-1.00920853E+02+4.86648027E+00+6.45174583E-02-2.45246679E-05    3
-1.77081536E-09+2.18648284E-12-3.20963786E+04+1.35846460E+01+0.00000000E+00    4
C7KET42O                C   7H  13O   2    0G   300.000  5000.000 1370.000    61
+2.56884614E+01+2.80095890E-02-9.25680532E-06+1.40530115E-09-8.03019698E-14    2
-4.20976441E+04-1.02650105E+02+4.70018599E+00+6.81280965E-02-3.21429326E-05    3
+3.33860657E-09+1.05751924E-12-3.41777201E+04+1.27950943E+01+0.00000000E+00    4
C7KET43O                C   7H  13O   2    0G   300.000  5000.000 1387.000    61
+2.52474702E+01+3.00387223E-02-1.02980700E-05+1.60151220E-09-9.30327317E-14    2
-4.15079135E+04-9.99196024E+01+4.22370120E+00+7.02977244E-02-3.51511137E-05    3
+5.96766285E-09+2.70620719E-13-3.33805928E+04+1.60319393E+01+0.00000000E+00    4
C7Y24                   C   7H  12O   2    0G   300.000  5000.000 1426.000    61
+2.33334638E+01+2.76457299E-02-9.17529929E-06+1.39740619E-09-8.00448780E-14    2
-6.12241187E+04-8.97827704E+01+4.39764101E+00+6.01180975E-02-2.22844519E-05    3
-1.91774372E-09+2.07240091E-12-5.36778370E+04+1.57433051E+01+0.00000000E+00    4
C7Y13                   C   7H  12O   2    0G   300.000  5000.000 1447.000    61
+2.43257239E+01+2.76226853E-02-9.33608747E-06+1.43914433E-09-8.31206829E-14    2
-5.80087604E+04-9.57614814E+01+3.61453518E+00+6.43014140E-02-2.64063505E-05    3
-1.08740222E-10+1.75733289E-12-4.98378626E+04+1.93018610E+01+0.00000000E+00    4
C7Y35                   C   7H  12O   2    0G   300.000  5000.000 1471.000    61
+2.29699639E+01+2.87451681E-02-9.71038176E-06+1.49572805E-09-8.63256686E-14    2
-6.08462735E+04-8.87044158E+01+3.89935666E+00+6.19920452E-02-2.45872500E-05    3
-3.61187603E-10+1.67912831E-12-5.32377873E+04+1.74838991E+01+0.00000000E+00    4
C7H14OOH1-2O            C   7H  15O   3    0G   300.000  5000.000 1684.000    81
+2.86766807E+01+3.64408431E-02-1.31971670E-05+2.13690883E-09-1.27860944E-13    2
-3.90828265E+04-1.15502906E+02+1.33099069E+00+9.67180192E-02-5.95878979E-05    3
+1.67058984E-08-1.64229299E-12-2.98431017E+04+3.17711823E+01+0.00000000E+00    4
C7H14OOH1-3O            C   7H  15O   3    0G   300.000  5000.000 1684.000    81
+2.86766807E+01+3.64408431E-02-1.31971670E-05+2.13690883E-09-1.27860944E-13    2
-3.90828265E+04-1.15502906E+02+1.33099069E+00+9.67180192E-02-5.95878979E-05    3
+1.67058984E-08-1.64229299E-12-2.98431017E+04+3.17711823E+01+0.00000000E+00    4
C7H14OOH1-4O            C   7H  15O   3    0G   300.000  5000.000 1684.000    81
+2.86766807E+01+3.64408431E-02-1.31971670E-05+2.13690883E-09-1.27860944E-13    2
-3.90828265E+04-1.15502906E+02+1.33099069E+00+9.67180192E-02-5.95878979E-05    3
+1.67058984E-08-1.64229299E-12-2.98431017E+04+3.17711823E+01+0.00000000E+00    4
C7H14OOH1-5O            C   7H  15O   3    0G   300.000  5000.000 1684.000    81
+2.86766807E+01+3.64408431E-02-1.31971670E-05+2.13690883E-09-1.27860944E-13    2
-3.90828265E+04-1.15502906E+02+1.33099069E+00+9.67180192E-02-5.95878979E-05    3
+1.67058984E-08-1.64229299E-12-2.98431017E+04+3.17711823E+01+0.00000000E+00    4
C7H14OOH2-1O            C   7H  15O   3    0G   300.000  5000.000 1407.000    81
+3.01497835E+01+3.22726460E-02-1.09797155E-05+1.69856254E-09-9.83026609E-14    2
-3.95955853E+04-1.23037063E+02+3.08548854E+00+9.51206736E-02-6.59996503E-05    3
+2.32444319E-08-3.27657401E-12-3.02456778E+04+2.23002772E+01+0.00000000E+00    4
C7H14OOH2-3O            C   7H  15O   3    0G   300.000  5000.000 1413.000    81
+3.02806950E+01+3.17579006E-02-1.07133963E-05+1.64778485E-09-9.49745325E-14    2
-4.14328088E+04-1.24204145E+02+3.01287651E+00+9.81864399E-02-7.25210341E-05    3
+2.76884286E-08-4.27353522E-12-3.23391710E+04+2.10962805E+01+0.00000000E+00    4
C7H14OOH2-4O            C   7H  15O   3    0G   300.000  5000.000 1413.000    81
+3.02806950E+01+3.17579006E-02-1.07133963E-05+1.64778485E-09-9.49745325E-14    2
-4.14328088E+04-1.24204145E+02+3.01287651E+00+9.81864399E-02-7.25210341E-05    3
+2.76884286E-08-4.27353522E-12-3.23391710E+04+2.10962805E+01+0.00000000E+00    4
C7H14OOH2-5O            C   7H  15O   3    0G   300.000  5000.000 1413.000    81
+3.02806950E+01+3.17579006E-02-1.07133963E-05+1.64778485E-09-9.49745325E-14    2
-4.14328088E+04-1.24204145E+02+3.01287651E+00+9.81864399E-02-7.25210341E-05    3
+2.76884286E-08-4.27353522E-12-3.23391710E+04+2.10962805E+01+0.00000000E+00    4
C7H14OOH2-6O            C   7H  15O   3    0G   300.000  5000.000 1413.000    81
+3.02806950E+01+3.17579006E-02-1.07133963E-05+1.64778485E-09-9.49745325E-14    2
-4.14328088E+04-1.24204145E+02+3.01287651E+00+9.81864399E-02-7.25210341E-05    3
+2.76884286E-08-4.27353522E-12-3.23391710E+04+2.10962805E+01+0.00000000E+00    4
C7H14OOH3-1O            C   7H  15O   3    0G   300.000  5000.000 1407.000    81
+3.01497835E+01+3.22726460E-02-1.09797155E-05+1.69856254E-09-9.83026609E-14    2
-3.95955853E+04-1.23037063E+02+3.08548854E+00+9.51206736E-02-6.59996503E-05    3
+2.32444319E-08-3.27657401E-12-3.02456778E+04+2.23002772E+01+0.00000000E+00    4
C7H14OOH3-2O            C   7H  15O   3    0G   300.000  5000.000 1413.000    81
+3.02806950E+01+3.17579006E-02-1.07133963E-05+1.64778485E-09-9.49745325E-14    2
-4.14328088E+04-1.24204145E+02+3.01287651E+00+9.81864399E-02-7.25210341E-05    3
+2.76884286E-08-4.27353522E-12-3.23391710E+04+2.10962805E+01+0.00000000E+00    4
C7H14OOH3-4O            C   7H  15O   3    0G   300.000  5000.000 1413.000    81
+3.02806950E+01+3.17579006E-02-1.07133963E-05+1.64778485E-09-9.49745325E-14    2
-4.14328088E+04-1.24204145E+02+3.01287651E+00+9.81864399E-02-7.25210341E-05    3
+2.76884286E-08-4.27353522E-12-3.23391710E+04+2.10962805E+01+0.00000000E+00    4
C7H14OOH3-5O            C   7H  15O   3    0G   300.000  5000.000 1413.000    81
+3.02806950E+01+3.17579006E-02-1.07133963E-05+1.64778485E-09-9.49745325E-14    2
-4.14328088E+04-1.24204145E+02+3.01287651E+00+9.81864399E-02-7.25210341E-05    3
+2.76884286E-08-4.27353522E-12-3.23391710E+04+2.10962805E+01+0.00000000E+00    4
C7H14OOH3-6O            C   7H  15O   3    0G   300.000  5000.000 1413.000    81
+3.02806950E+01+3.17579006E-02-1.07133963E-05+1.64778485E-09-9.49745325E-14    2
-4.14328088E+04-1.24204145E+02+3.01287651E+00+9.81864399E-02-7.25210341E-05    3
+2.76884286E-08-4.27353522E-12-3.23391710E+04+2.10962805E+01+0.00000000E+00    4
C7H14OOH3-7O            C   7H  15O   3    0G   300.000  5000.000 1407.000    81
+3.01497835E+01+3.22726460E-02-1.09797155E-05+1.69856254E-09-9.83026609E-14    2
-3.95955853E+04-1.23037063E+02+3.08548854E+00+9.51206736E-02-6.59996503E-05    3
+2.32444319E-08-3.27657401E-12-3.02456778E+04+2.23002772E+01+0.00000000E+00    4
C7H14OOH4-1O            C   7H  15O   3    0G   300.000  5000.000 1407.000    81
+3.01497835E+01+3.22726460E-02-1.09797155E-05+1.69856254E-09-9.83026609E-14    2
-3.95955853E+04-1.23037063E+02+3.08548854E+00+9.51206736E-02-6.59996503E-05    3
+2.32444319E-08-3.27657401E-12-3.02456778E+04+2.23002772E+01+0.00000000E+00    4
C7H14OOH4-2O            C   7H  15O   3    0G   300.000  5000.000 1413.000    81
+3.02806950E+01+3.17579006E-02-1.07133963E-05+1.64778485E-09-9.49745325E-14    2
-4.14328088E+04-1.24204145E+02+3.01287651E+00+9.81864399E-02-7.25210341E-05    3
+2.76884286E-08-4.27353522E-12-3.23391710E+04+2.10962805E+01+0.00000000E+00    4
C7H14OOH4-3O            C   7H  15O   3    0G   300.000  5000.000 1413.000    81
+3.02806950E+01+3.17579006E-02-1.07133963E-05+1.64778485E-09-9.49745325E-14    2
-4.14328088E+04-1.24204145E+02+3.01287651E+00+9.81864399E-02-7.25210341E-05    3
+2.76884286E-08-4.27353522E-12-3.23391710E+04+2.10962805E+01+0.00000000E+00    4
C6H11O13-6              C   6H  11O   1    0G   300.000  5000.000 1412.000    31
+1.94680493E+01+2.55210612E-02-8.62688975E-06+1.32887037E-09-7.66797753E-14    2
-4.82503956E+03-7.66455390E+01-8.55042113E+00+9.93712909E-02-8.38485087E-05    3
+3.62206697E-08-6.24312731E-12+3.95319530E+03+7.06614274E+01+0.00000000E+00    4
C6H11O14-6              C   6H  11O   1    0G   300.000  5000.000 1455.000    21
+1.82831468E+01+2.54265745E-02-8.27252851E-06+1.24123104E-09-7.03046026E-14    2
-1.42244253E+04-7.02944830E+01-7.80524702E+00+9.37481232E-02-7.60016637E-05    3
+3.12611899E-08-5.06939758E-12-6.15964922E+03+6.67633621E+01+0.00000000E+00    4
C6H11O15-6              C   6H  11O   1    0G   300.000  5000.000 1444.000    11
+1.87856469E+01+2.59182642E-02-8.54662736E-06+1.29454658E-09-7.38246342E-14    2
-1.67718783E+04-7.84622939E+01-8.38439662E+00+9.57209767E-02-7.64661564E-05    3
+3.08782447E-08-4.92187508E-12-8.21380764E+03+6.47980999E+01+0.00000000E+00    4
C6H11O23-1              C   6H  11O   1    0G   300.000  5000.000 1428.000    41
+2.09510264E+01+2.32219824E-02-7.70555586E-06+1.17228694E-09-6.70636135E-14    2
-6.04704320E+03-8.35825137E+01-4.92079122E+00+9.07221617E-02-7.48659944E-05    3
+3.12724603E-08-5.16926400E-12+2.03286829E+03+5.25244419E+01+0.00000000E+00    4
C6H11O23-6              C   6H  11O   1    0G   300.000  5000.000 1428.000    41
+2.09510264E+01+2.32219824E-02-7.70555586E-06+1.17228694E-09-6.70636135E-14    2
-6.04704320E+03-8.35825137E+01-4.92079122E+00+9.07221617E-02-7.48659944E-05    3
+3.12724603E-08-5.16926400E-12+2.03286829E+03+5.25244419E+01+0.00000000E+00    4
C6H11O24-1              C   6H  11O   1    0G   300.000  5000.000 1418.000    31
+1.97676292E+01+2.48505263E-02-8.30594789E-06+1.26961939E-09-7.28648539E-14    2
-6.74869207E+03-7.88109458E+01-8.34495598E+00+1.01028943E-01-8.78699575E-05    3
+3.89477222E-08-6.83884937E-12+1.82049644E+03+6.82011830E+01+0.00000000E+00    4
C6H11O24-6              C   6H  11O   1    0G   300.000  5000.000 1418.000    31
+1.97676292E+01+2.48505263E-02-8.30594789E-06+1.26961939E-09-7.28648539E-14    2
-6.74869207E+03-7.88109458E+01-8.34495598E+00+1.01028943E-01-8.78699575E-05    3
+3.89477222E-08-6.83884937E-12+1.82049644E+03+6.82011830E+01+0.00000000E+00    4
C6H11O34-1              C   6H  11O   1    0G   300.000  5000.000 1428.000    41
+2.09510264E+01+2.32219824E-02-7.70555586E-06+1.17228694E-09-6.70636135E-14    2
-6.04704320E+03-8.35825137E+01-4.92079122E+00+9.07221617E-02-7.48659944E-05    3
+3.12724603E-08-5.16926400E-12+2.03286829E+03+5.25244419E+01+0.00000000E+00    4
C6Y2-1J                 C   6H  11O   1    0G   300.000  5000.000 1396.000    51
+2.04383273E+01+2.38253206E-02-8.04100895E-06+1.23762461E-09-7.13843846E-14    2
-2.16182253E+04-7.85923730E+01+1.75975194E+00+6.42520985E-02-3.96352767E-05    3
+1.15685286E-08-1.20137340E-12-1.48945661E+04+2.27202794E+01+0.00000000E+00    4
C6Y3-6J                 C   6H  11O   1    0G   300.000  5000.000 1428.000    51
+1.93145300E+01+2.40496101E-02-7.97552707E-06+1.21393244E-09-6.95022464E-14    2
-1.87180946E+04-7.10938989E+01+3.01181403E+00+5.23666148E-02-2.00629431E-05    3
-1.05670148E-09+1.64429373E-12-1.22517682E+04+1.96394582E+01+0.00000000E+00    4
C6Y3-1J                 C   6H  11O   1    0G   300.000  5000.000 1428.000    51
+1.93145300E+01+2.40496101E-02-7.97552707E-06+1.21393244E-09-6.95022464E-14    2
-1.87180946E+04-7.10938989E+01+3.01181403E+00+5.23666148E-02-2.00629431E-05    3
-1.05670148E-09+1.64429373E-12-1.22517682E+04+1.96394582E+01+0.00000000E+00    4
C7H14-1                 C   7H  14    0    0G   300.000  5000.000 1392.000    51
+2.10516278E+01+3.12760197E-02-1.06771829E-05+1.65550145E-09-9.59594932E-14    2
-1.83777234E+04-8.41750939E+01-8.09358679E-01+7.89648824E-02-4.95897128E-05    3
+1.57930253E-08-2.02821634E-12-1.04146627E+04+3.44853698E+01+0.00000000E+00    4
C7H14-2                 C   7H  14    0    0G   300.000  5000.000 1389.000    51
+2.06209791E+01+3.15553139E-02-1.07554876E-05+1.66593057E-09-9.64967953E-14    2
-1.95694445E+04-8.23986766E+01-5.38953650E-02+7.44295393E-02-4.28542682E-05    3
+1.17521061E-08-1.16517055E-12-1.18188874E+04+3.06085980E+01+0.00000000E+00    4
C7H14-3                 C   7H  14    0    0G   300.000  5000.000 1388.000    51
+2.03621010E+01+3.16779587E-02-1.07777153E-05+1.66742019E-09-9.65068542E-14    2
-1.94856293E+04-8.10623354E+01-4.98371307E-01+7.49068336E-02-4.30333630E-05    3
+1.17133021E-08-1.13719824E-12-1.16707063E+04+3.29566580E+01+0.00000000E+00    4
C7H131-3                C   7H  13    0    0G   300.000  5000.000 1384.000    41
+2.14156908E+01+2.85177236E-02-9.66514723E-06+1.49210849E-09-8.62535195E-14    2
-1.70979838E+03-8.60030226E+01-5.60862522E-01+7.54326016E-02-4.60711095E-05    3
+1.34950109E-08-1.45966663E-12+6.32990830E+03+3.35375654E+01+0.00000000E+00    4
C7H131-4                C   7H  13    0    0G   300.000  5000.000 1393.000    51
+1.95903002E+01+2.99096858E-02-1.01928469E-05+1.57855426E-09-9.14249512E-14    2
+5.42884260E+03-7.29326843E+01+7.59883219E-01+6.65218933E-02-3.38705045E-05    3
+6.62244871E-09-5.39889345E-14+1.26842125E+04+3.07767256E+01+0.00000000E+00    4
C7H131-5                C   7H  13    0    0G   300.000  5000.000 1393.000    51
+1.95903002E+01+2.99096858E-02-1.01928469E-05+1.57855426E-09-9.14249512E-14    2
+5.42884260E+03-7.29326843E+01+7.59883219E-01+6.65218933E-02-3.38705045E-05    3
+6.62244871E-09-5.39889345E-14+1.26842125E+04+3.07767256E+01+0.00000000E+00    4
C7H131-6                C   7H  13    0    0G   300.000  5000.000 1393.000    51
+1.95903002E+01+2.99096858E-02-1.01928469E-05+1.57855426E-09-9.14249512E-14    2
+5.42884260E+03-7.29326843E+01+7.59883219E-01+6.65218933E-02-3.38705045E-05    3
+6.62244871E-09-5.39889345E-14+1.26842125E+04+3.07767256E+01+0.00000000E+00    4
C7H131-7                C   7H  13    0    0G   300.000  5000.000 1393.000    51
+2.04254451E+01+2.93645160E-02-1.00400399E-05+1.55828940E-09-9.03875243E-14    2
+6.75757861E+03-7.80202543E+01-4.40736730E-01+7.55083258E-02-4.85768313E-05    3
+1.60730287E-08-2.17974149E-12+1.43050908E+04+3.50343173E+01+0.00000000E+00    4
C7H132-4                C   7H  13    0    0G   300.000  5000.000 1389.000    41
+2.02204603E+01+2.98619421E-02-1.01919239E-05+1.58015892E-09-9.15931884E-14    2
-2.52466923E+03-8.14726926E+01-3.72763979E-01+7.27705155E-02-4.24262213E-05    3
+1.17101335E-08-1.15624520E-12+5.15547887E+03+3.09838851E+01+0.00000000E+00    4
C7H132-5                C   7H  13    0    0G   300.000  5000.000 1391.000    51
+1.90854765E+01+3.01791168E-02-1.02513232E-05+1.58415277E-09-9.16099642E-14    2
+4.31614862E+03-7.06165152E+01+1.82382661E+00+6.10673441E-02-2.62220491E-05    3
+2.14472121E-09+8.93751848E-13+1.12216271E+04+2.53795314E+01+0.00000000E+00    4
C7H132-6                C   7H  13    0    0G   300.000  5000.000 1391.000    51
+1.90854765E+01+3.01791168E-02-1.02513232E-05+1.58415277E-09-9.16099642E-14    2
+4.31614862E+03-7.06165152E+01+1.82382661E+00+6.10673441E-02-2.62220491E-05    3
+2.14472121E-09+8.93751848E-13+1.12216271E+04+2.53795314E+01+0.00000000E+00    4
C7H132-7                C   7H  13    0    0G   300.000  5000.000 1390.000    51
+1.99821175E+01+2.96591221E-02-1.01244293E-05+1.56973641E-09-9.09863758E-14    2
+5.57188959E+03-7.61641862E+01+3.58569522E-01+7.07856603E-02-4.15780734E-05    3
+1.18775321E-08-1.28395050E-12+1.28940839E+04+3.09582265E+01+0.00000000E+00    4
C7H133-1                C   7H  13    0    0G   300.000  5000.000 1389.000    51
+1.97137107E+01+2.97943652E-02-1.01517896E-05+1.57209319E-09-9.10491100E-14    2
+5.66002000E+03-7.47727706E+01-7.85839985E-02+7.12349539E-02-4.17259682E-05    3
+1.18251338E-08-1.25384179E-12+1.30410765E+04+3.32716438E+01+0.00000000E+00    4
C7H133-5                C   7H  13    0    0G   300.000  5000.000 1388.000    41
+1.99813268E+01+2.99618307E-02-1.02051724E-05+1.58014428E-09-9.15119629E-14    2
-2.44655429E+03-8.02443024E+01-8.13432333E-01+7.32810249E-02-4.26690697E-05    3
+1.17112103E-08-1.13686121E-12+5.30153685E+03+3.33028462E+01+0.00000000E+00    4
C7H133-6                C   7H  13    0    0G   300.000  5000.000 1388.000    51
+1.88327779E+01+3.03047716E-02-1.02765174E-05+1.58631403E-09-9.16678097E-14    2
+4.39301285E+03-6.93248547E+01+1.39520323E+00+6.14606183E-02-2.62663084E-05    3
+2.02811054E-09+9.36702991E-13+1.13677716E+04+2.76569852E+01+0.00000000E+00    4
C7H133-7                C   7H  13    0    0G   300.000  5000.000 1389.000    51
+1.97137107E+01+2.97943652E-02-1.01517896E-05+1.57209319E-09-9.10491100E-14    2
+5.66002000E+03-7.47727706E+01-7.85839985E-02+7.12349539E-02-4.17259682E-05    3
+1.18251338E-08-1.25384179E-12+1.30410765E+04+3.32716438E+01+0.00000000E+00    4
C7H13-1D3O              C   7H  13O   1    0G   300.000  5000.000 1385.000    51
+2.45962638E+01+2.91695918E-02-1.01515243E-05+1.59445051E-09-9.32566850E-14    2
-1.27137607E+04-9.96395968E+01+1.75836665E+00+7.85031672E-02-5.03690559E-05    3
+1.64406880E-08-2.20903728E-12-4.28436460E+03+2.46022100E+01+0.00000000E+00    4
C7H13-2D4O              C   7H  13O   1    0G   300.000  5000.000 1383.000    51
+2.41090151E+01+2.95611974E-02-1.02814801E-05+1.61418484E-09-9.43829333E-14    2
-1.38756865E+04-9.75312193E+01+2.63531821E+00+7.36578610E-02-4.33517009E-05    3
+1.23129314E-08-1.34071479E-12-5.71335565E+03+2.01138895E+01+0.00000000E+00    4
C7H13-3D5O              C   7H  13O   1    0G   300.000  5000.000 1383.000    51
+2.37587144E+01+2.98416387E-02-1.03744412E-05+1.62830253E-09-9.51890868E-14    2
-1.37728890E+04-9.57179560E+01+2.19575759E+00+7.38969654E-02-4.30597626E-05    3
+1.19763351E-08-1.24916735E-12-5.55965639E+03+2.24865296E+01+0.00000000E+00    4
C7H14OH-1J2             C   7H  15O   1    0G   300.000  5000.000 1396.000    71
+2.38166116E+01+3.29487814E-02-1.12036524E-05+1.73236311E-09-1.00218147E-13    2
-2.87703608E+04-9.19434776E+01+1.21072127E+00+8.32765482E-02-5.34939093E-05    3
+1.77237371E-08-2.40178894E-12-2.06442678E+04+3.03879690E+01+0.00000000E+00    4
C7H14OH-2J1             C   7H  15O   1    0G   300.000  5000.000 1402.000    71
+2.50087998E+01+3.15305124E-02-1.06261019E-05+1.63312194E-09-9.40751455E-14    2
-2.97161468E+04-9.92807674E+01+8.16287767E-01+9.08578310E-02-6.71105637E-05    3
+2.63947068E-08-4.28593595E-12-2.15950059E+04+2.96490882E+01+0.00000000E+00    4
C7H14OH-2J3             C   7H  15O   1    0G   300.000  5000.000 1401.000    71
+2.41756177E+01+3.20133170E-02-1.07458095E-05+1.64715331E-09-9.47106929E-14    2
-3.06787328E+04-9.43545895E+01+9.10348667E-01+8.72019493E-02-6.09956660E-05    3
+2.25368413E-08-3.43473439E-12-2.27001132E+04+3.02657448E+01+0.00000000E+00    4
C7H14OH-3J2             C   7H  15O   1    0G   300.000  5000.000 1401.000    71
+2.41756177E+01+3.20133170E-02-1.07458095E-05+1.64715331E-09-9.47106929E-14    2
-3.06787328E+04-9.43545895E+01+9.10348667E-01+8.72019493E-02-6.09956660E-05    3
+2.25368413E-08-3.43473439E-12-2.27001132E+04+3.02657448E+01+0.00000000E+00    4
C7H14OH-3J4             C   7H  15O   1    0G   300.000  5000.000 1401.000    71
+2.41756177E+01+3.20133170E-02-1.07458095E-05+1.64715331E-09-9.47106929E-14    2
-3.06787328E+04-9.43545895E+01+9.10348667E-01+8.72019493E-02-6.09956660E-05    3
+2.25368413E-08-3.43473439E-12-2.27001132E+04+3.02657448E+01+0.00000000E+00    4
C7H14OH-4J3             C   7H  15O   1    0G   300.000  5000.000 1401.000    71
+2.41756177E+01+3.20133170E-02-1.07458095E-05+1.64715331E-09-9.47106929E-14    2
-3.06787328E+04-9.43545895E+01+9.10348667E-01+8.72019493E-02-6.09956660E-05    3
+2.25368413E-08-3.43473439E-12-2.27001132E+04+3.02657448E+01+0.00000000E+00    4
C7H14OH-1O2-2           C   7H  15O   3    0G   300.000  5000.000 1403.000    81
+2.96517284E+01+3.27070176E-02-1.11327901E-05+1.72285104E-09-9.97346708E-14    2
-4.94593269E+04-1.19933256E+02+8.62497819E-01+1.01693666E-01-7.43995933E-05    3
+2.81050374E-08-4.31255025E-12-3.96992260E+04+3.39577229E+01+0.00000000E+00    4
C7H14OH-2O2-1           C   7H  15O   3    0G   300.000  5000.000 1401.000    81
+2.87755285E+01+3.34750290E-02-1.14005874E-05+1.76476211E-09-1.02173530E-13    2
-4.91233276E+04-1.14722340E+02+5.37268604E-01+1.02515862E-01-7.68815510E-05    3
+3.03521838E-08-4.92329087E-12-3.96260600E+04+3.58384566E+01+0.00000000E+00    4
C7H14OH-2O2-3           C   7H  15O   3    0G   300.000  5000.000 1407.000    81
+2.91474754E+01+3.26332166E-02-1.09950902E-05+1.68957012E-09-9.73167191E-14    2
-5.09733381E+04-1.17279245E+02+9.53439399E-01+1.04452051E-01-8.20570973E-05    3
+3.39454494E-08-5.71650860E-12-4.18203504E+04+3.19524737E+01+0.00000000E+00    4
C7H14OH-3O2-2           C   7H  15O   3    0G   300.000  5000.000 1407.000    81
+2.91474754E+01+3.26332166E-02-1.09950902E-05+1.68957012E-09-9.73167191E-14    2
-5.09733381E+04-1.17279245E+02+9.53439399E-01+1.04452051E-01-8.20570973E-05    3
+3.39454494E-08-5.71650860E-12-4.18203504E+04+3.19524737E+01+0.00000000E+00    4
C7H14OH-3O2-4           C   7H  15O   3    0G   300.000  5000.000 1407.000    81
+2.91474754E+01+3.26332166E-02-1.09950902E-05+1.68957012E-09-9.73167191E-14    2
-5.09733381E+04-1.17279245E+02+9.53439399E-01+1.04452051E-01-8.20570973E-05    3
+3.39454494E-08-5.71650860E-12-4.18203504E+04+3.19524737E+01+0.00000000E+00    4
C7H14OH-4O2-3           C   7H  15O   3    0G   300.000  5000.000 1407.000    81
+2.91474754E+01+3.26332166E-02-1.09950902E-05+1.68957012E-09-9.73167191E-14    2
-5.09733381E+04-1.17279245E+02+9.53439399E-01+1.04452051E-01-8.20570973E-05    3
+3.39454494E-08-5.71650860E-12-4.18203504E+04+3.19524737E+01+0.00000000E+00    4
C5D2Y1-1R               C   5H   7O   1    0G   300.000  5000.000 1390.000    31
+1.58396423E+01+1.66571765E-02-5.74155776E-06+8.96152306E-10-5.21898413E-14    2
-5.43955462E+03-5.57243534E+01+7.67163837E-01+5.23888982E-02-3.85650887E-05    3
+1.48263722E-08-2.35263797E-12-2.36668558E+02+2.50746199E+01+0.00000000E+00    4
C3Y1-3OR                C   3H   5O   2    0G   300.000  5000.000 1409.000    31
+1.24458641E+01+1.15135588E-02-3.89008277E-06+5.99667928E-10-3.46406544E-14    2
-2.78997305E+04-3.52984011E+01+2.64167269E+00+2.94283641E-02-1.29127845E-05    3
+3.88757872E-10+7.42968763E-13-2.41114860E+04+1.89330066E+01+0.00000000E+00    4
C4Y1-3OR                C   4H   7O   2    0G   300.000  5000.000 1417.000    31
+1.64998473E+01+1.58390093E-02-5.41015815E-06+8.39905247E-10-4.87505919E-14    2
-2.64232542E+04-5.83737300E+01+3.94683511E+00+3.65984570E-02-1.24268392E-05    3
-2.56058969E-09+1.66288190E-12-2.13506683E+04+1.18427218E+01+0.00000000E+00    4
C6D2Y1                  C   6H  10O   1    0G   300.000  5000.000 1392.000    41
+1.95305471E+01+2.32320952E-02-7.99721990E-06+1.24699364E-09-7.25687500E-14    2
-2.85719761E+04-7.57135584E+01-2.69585026E-01+6.98099901E-02-5.04217305E-05    3
+1.90982509E-08-2.99716926E-12-2.16923258E+04+3.05709242E+01+0.00000000E+00    4
C6D2Y1-1R               C   6H   9O   1    0G   300.000  5000.000 1392.000    41
+1.91108039E+01+2.11064142E-02-7.27838190E-06+1.13627682E-09-6.61818880E-14    2
-9.60886866E+03-7.17888495E+01+5.03660007E-01+6.50190464E-02-4.73912739E-05    3
+1.80513164E-08-2.84079598E-12-3.16399550E+03+2.80316159E+01+0.00000000E+00    4
H15DE25DM               C   8H  14    0    0G   300.000  5000.000 1395.000    51
+2.25355644E+01+3.23955734E-02-1.10270814E-05+1.70640907E-09-9.87758061E-14    2
-1.04808866E+04-9.19784905E+01-1.71853441E+00+8.82613783E-02-6.03140500E-05    3
+2.15862289E-08-3.19690882E-12-1.95255748E+03+3.86048681E+01+0.00000000E+00    4
H15DE25DM-S             C   8H  13    0    0G   300.000  5000.000 1395.000    41
+2.21422958E+01+3.06966055E-02-1.04617380E-05+1.62037747E-09-9.38578511E-14    2
+6.56045671E+03-9.04059585E+01-2.04235551E+00+8.66261688E-02-5.99110976E-05    3
+2.15551630E-08-3.18976697E-12+1.50224279E+04+3.96917763E+01+0.00000000E+00    4
H15DE25DM-A             C   8H  13    0    0G   300.000  5000.000 1391.000    41
+2.33282646E+01+2.93694154E-02-9.94258906E-06+1.53368063E-09-8.86030202E-14    2
+7.37319036E+03-9.55902415E+01-2.21863377E+00+8.91652629E-02-6.33360636E-05    3
+2.32007379E-08-3.46329567E-12+1.61971179E+04+4.15116620E+01+0.00000000E+00    4
H15DE25DM-AO            C   8H  13O   1    0G   300.000  5000.000 1378.000    51
+2.50985951E+01+3.15085628E-02-1.10076915E-05+1.73332426E-09-1.01557468E-13    2
-2.49465338E+03-1.01097942E+02+3.03691957E+00+7.50640438E-02-4.17779534E-05    3
+1.07915725E-08-9.97734397E-13+6.11649780E+03+2.04746031E+01+0.00000000E+00    4
H15DE25DM-SO            C   8H  13O   1    0G   300.000  5000.000 1388.000    51
+2.60152179E+01+3.04295766E-02-1.05676513E-05+1.65746547E-09-9.68470091E-14    2
-4.79568520E+03-1.06442472E+02+9.30464015E-01+8.71669873E-02-5.99582593E-05    3
+2.15026041E-08-3.21687573E-12+4.19310073E+03+2.90924508E+01+0.00000000E+00    4
H15DE2M-T               C   7H  11    0    0G   300.000  5000.000 1389.000    41
+1.90144729E+01+2.61932198E-02-9.01183878E-06+1.40455988E-09-8.17075251E-14    2
+2.35551101E+04-7.15568628E+01+3.88856066E-01+6.70215700E-02-4.29671268E-05    3
+1.42489875E-08-1.96105571E-12+3.03627273E+04+2.95444186E+01+0.00000000E+00    4
IC4H7CHO                C   5H   8O   1    0G   300.000  5000.000 1391.000    31
+1.59171638E+01+1.93357284E-02-6.70857943E-06+1.05155191E-09-6.14175906E-14    2
-2.16140735E+04-5.67616631E+01-1.20982776E+00+5.92603375E-02-4.26960089E-05    3
+1.60356164E-08-2.49347521E-12-1.56205327E+04+3.53137305E+01+0.00000000E+00    4
C8H141-5,3-4            C   8H  14    0    0G   300.000  5000.000 1396.000    51
+2.30690680E+01+3.23154042E-02-1.10795683E-05+1.72276354E-09-1.00052582E-13    2
-8.91240214E+03-9.49655754E+01-2.52713194E+00+9.28837673E-02-6.67176819E-05    3
+2.53683579E-08-4.01212661E-12-4.55965940E+01+4.23180878E+01+0.00000000E+00    4
C8H131-5,3-4,TA         C   8H  13    0    0G   300.000  5000.000 1394.000    41
+2.22822575E+01+3.10651867E-02-1.06940907E-05+1.66739777E-09-9.70243450E-14    2
+7.57680613E+03-9.19858764E+01-3.23996819E+00+9.13494930E-02-6.60037456E-05    3
+2.51706078E-08-3.99030974E-12+1.64345368E+04+4.49498860E+01+0.00000000E+00    4
C6H101-3,3              C   6H  10    0    0G   300.000  5000.000 1395.000    31
+1.69678361E+01+2.28868236E-02-7.78758381E-06+1.20465198E-09-6.97080856E-14    2
-2.97276905E+03-6.58632941E+01-3.01310455E-02+6.43105079E-02-4.75083462E-05    3
+1.89877768E-08-3.17681035E-12+2.82367411E+03+2.49254708E+01+0.00000000E+00    4
C8H131-5,3-4,TAO        C   8H  13O   1    0G   300.000  5000.000 1394.000    51
+2.70579050E+01+2.84726632E-02-9.66434779E-06+1.49337149E-09-8.63788413E-14    2
-4.43111126E+03-1.12228392E+02+1.00679908E+00+8.90191278E-02-6.27963646E-05    3
+2.24161585E-08-3.20587060E-12+4.56422741E+03+2.76546640E+01+0.00000000E+00    4
C8H141-5,3  8/25/15     C   8H  14    0    0G   300.000  5000.000 1392.000    51
+2.25173982E+01+3.26748629E-02-1.11807923E-05+1.73629966E-09-1.00752481E-13    2
-8.96062790E+03-9.10857551E+01-1.02072126E+00+8.47808555E-02-5.47568199E-05    3
+1.81792070E-08-2.47335881E-12-4.53248586E+02+3.64247438E+01+0.00000000E+00    4
C8H131-5,3,TA           C   8H  13    0    0G   300.000  5000.000 1389.000    41
+2.16161787E+01+3.14326704E-02-1.07786324E-05+1.67632587E-09-9.73755313E-14    2
+7.60897211E+03-8.80384104E+01-5.03201172E-01+7.78854227E-02-4.63156182E-05    3
+1.32834166E-08-1.42623050E-12+1.58388712E+04+3.26514434E+01+0.00000000E+00    4
C8H131-5,3,SA           C   8H  13    0    0G   300.000  5000.000 1392.000    41
+2.21141889E+01+3.09871348E-02-1.06198459E-05+1.65100088E-09-9.58788408E-14    2
+8.08509780E+03-9.01448021E+01-1.32185914E+00+8.30473789E-02-5.42213233E-05    3
+1.80737386E-08-2.45105483E-12+1.65183103E+04+3.67169651E+01+0.00000000E+00    4
C8H131-5,3,PA           C   8H  13    0    0G   300.000  5000.000 1389.000    41
+2.32085707E+01+2.97529224E-02-1.01333635E-05+1.56925634E-09-9.09001242E-14    2
+8.95338901E+03-9.40777602E+01-1.57063382E+00+8.60080913E-02-5.83884368E-05    3
+2.02048105E-08-2.83115953E-12+1.77015232E+04+3.95476224E+01+0.00000000E+00    4
C8H131-5,3,TAO          C   8H  13O   1    0G   300.000  5000.000 1396.000    51
+2.16638860E+01+2.77253448E-02-9.69375951E-06+1.67582120E-09-1.08059396E-13    2
-5.70300683E+03-9.33237797E+01+1.46771925E+00+7.67800622E-02-5.63189881E-05    3
+2.22689786E-08-3.64813515E-12+1.17475936E+03+1.45619856E+01+0.00000000E+00    4
C8H131-5,3,SAO          C   8H  13O   1    0G   300.000  5000.000 1385.000    51
+2.61023602E+01+3.05036647E-02-1.06268215E-05+1.67026867E-09-9.77389024E-14    2
-3.64744193E+03-1.06781316E+02+1.60953926E+00+8.39738786E-02-5.49469234E-05    3
+1.84255257E-08-2.56040058E-12+5.33713436E+03+2.62653941E+01+0.00000000E+00    4
C8H131-5,3,PAO          C   8H  13O   1    0G   300.000  5000.000 1374.000    51
+2.51902631E+01+3.15630048E-02-1.10568300E-05+1.74424175E-09-1.02327221E-13    2
-1.34401684E+03-1.01448477E+02+3.91532442E+00+7.10319966E-02-3.55623644E-05    3
+6.98595095E-09-1.83465840E-13+7.22911524E+03+1.67145758E+01+0.00000000E+00    4
C7H111-5,3,6P           C   7H  11    0    0G   300.000  5000.000 1396.000    41
+1.95787047E+01+2.54213538E-02-8.68127275E-06+1.34629701E-09-7.80464853E-14    2
+2.58537943E+04-7.44112330E+01-6.76848821E-01+7.38082653E-02-5.35945220E-05    3
+2.06293915E-08-3.29701110E-12+3.28160434E+04+3.40518079E+01+0.00000000E+00    4
C8H142-6   8/25/15      C   8H  14    0    0G   300.000  5000.000 1386.000    51
+2.20960852E+01+3.27887472E-02-1.11700037E-05+1.72970378E-09-1.00179059E-13    2
-9.04951881E+03-8.92942652E+01+3.43524821E-01+7.72359120E-02-4.34861460E-05    3
+1.12949093E-08-9.77995416E-13-8.37798357E+02+2.98241439E+01+0.00000000E+00    4
C8H132-6,SA             C   8H  13    0    0G   300.000  5000.000 1387.000    41
+2.16167233E+01+3.12260643E-02-1.06640216E-05+1.65409816E-09-9.59112187E-14    2
+8.03384556E+03-8.72194430E+01+2.20017932E-01+7.48621425E-02-4.21239973E-05    3
+1.07414215E-08-8.66560315E-13+1.61027987E+04+2.99517204E+01+0.00000000E+00    4
C8H132-6,PA             C   8H  13    0    0G   300.000  5000.000 1378.000    41
+2.29293875E+01+2.97187394E-02-1.00712335E-05+1.55505094E-09-8.99129602E-14    2
+8.77975921E+03-9.24517461E+01+1.05119796E-01+7.70150350E-02-4.48890925E-05    3
+1.19516688E-08-1.04377517E-12+1.72713386E+04+3.22058738E+01+0.00000000E+00    4
C8H132-6,SAO            C   8H  13O   1    0G   300.000  5000.000 1381.000    51
+2.54267504E+01+3.10421548E-02-1.08045689E-05+1.69716523E-09-9.92701997E-14    2
-3.28641768E+03-1.02872762E+02+3.34168622E+00+7.49917518E-02-4.18382842E-05    3
+1.06108028E-08-8.96488454E-13+5.24458399E+03+1.86128166E+01+0.00000000E+00    4
C8H132-6,PAO            C   8H  13O   1    0G   300.000  5000.000 2014.000    51
+1.99391776E+01+3.79081645E-02-1.37893231E-05+2.23770591E-09-1.34044177E-13    2
+1.42981257E+03-7.07923233E+01+6.30807632E+00+5.80374259E-02-1.75637726E-05    3
-2.70887760E-09+1.61702129E-12+7.07839485E+03+6.29344560E+00+0.00000000E+00    4
C7H111-5,1P             C   7H  11    0    0G   300.000  5000.000 1388.000    41
+1.91915682E+01+2.55013021E-02-8.65881522E-06+1.33796943E-09-7.73784878E-14    2
+2.60946287E+04-7.21387547E+01+8.16831855E-01+6.56745024E-02-4.14490949E-05    3
+1.32234876E-08-1.69289568E-12+3.27646149E+04+2.75442934E+01+0.00000000E+00    4
L-C6H4            H6W/94C   6H   4    0    0G   300.000  3000.00  1000.00      1
+1.27151820E+01+1.38396620E-02-4.37654400E-06+3.15416360E-10+4.66190260E-14    2
+5.70311480E+04-3.94646000E+01+2.95902250E-01+5.80533180E-02-6.77667560E-05    3
+4.33767620E-08-1.14188640E-11+6.00013710E+04+2.23189700E+01+0.00000000E+00    4
C-C6H4            H6W/94C   6H   4    0    0G   300.000  3000.00  1000.00      1
+1.38492090E+01+7.88079200E-03+1.82438360E-06-2.11691660E-09+3.74599770E-13    2
+4.74463400E+04-5.04049530E+01-3.09912680E+00+5.40305640E-02-4.08390040E-05    3
+1.07388370E-08+9.80784900E-13+5.22057110E+04+3.74152070E+01+0.00000000E+00    4
C6H3              H6W/94C   6H   3    0    0G   300.000  3000.00  1000.00      1
+5.81883430E+00+2.79334080E-02-1.78254270E-05+5.37025360E-09-6.17076270E-13    2
+8.51882500E+04-9.21478270E-01+1.17906190E+00+5.55473600E-02-7.30761680E-05    3
+5.20767360E-08-1.50469640E-11+8.56473120E+04+1.91791990E+01+0.00000000E+00    4
C6H2              P 1/93C   6H   2    0    0G   300.000  3000.00  1000.00      1
+1.32262810E+01+7.39043020E-03-2.27153810E-06+2.58752170E-10-5.53567410E-15    2
+8.05652580E+04-4.12011760E+01-1.59326240E+00+8.05301450E-02-1.48006490E-04    3
+1.33000310E-07-4.53323130E-11+8.32732270E+04+2.79808730E+01+0.00000000E+00    4
C6H6              G 6/01C   6H   6    0    0G   200.000  6000.000 1000.000     1
+1.10809576E+01+2.07176746E-02-7.52145991E-06+1.22320984E-09-7.36091279E-14    2
+4.30641035E+03-4.00413310E+01+5.04818632E-01+1.85020642E-02+7.38345881E-05    3
-1.18135741E-07+5.07210429E-11+8.55247913E+03+2.16412893E+01+9.96811598E+03    4
FULVENE                0C   6H   6    0    0G   200.000  5000.000 1000.00    0 1
+1.11035250E+01+2.06006850E-02-7.53022240E-06+1.23886950E-09-7.54159760E-14    2
+2.03618430E+04-3.66651970E+01-7.18131910E-01+3.79343120E-02+1.13988370E-05    3
-4.13335030E-08+1.80559270E-11+2.42238250E+04+2.78557140E+01+0.00000000E+00    4
C6H5              T04/02C   6H   5    0    0G   200.000  6000.000 1000.        1
+1.08444762E+01+1.73212473E-02-6.29233249E-06+1.02369961E-09-6.16216828E-14    2
+3.55598475E+04-3.53735134E+01+2.10306633E-01+2.04745507E-02+5.89743006E-05    3
-1.01534255E-07+4.47105660E-11+3.95468722E+04+2.52910455E+01+4.08610970E+04    4
C6H5OO     3/26/ 9 THERMC   6H   5O   2    0G   300.000  5000.000 1403.000    11
+1.67078262E+01+1.62326229E-02-5.47969630E-06+8.43510060E-10-4.86562431E-14    2
+8.14242915E+03-6.08346973E+01-2.99164672E+00+7.03857150E-02-6.34400574E-05    3
+2.91548920E-08-5.30706938E-12+1.41320240E+04+4.20142955E+01+0.00000000E+00    4
C6H5OOH    3/26/ 9 THERMC   6H   6O   2    0G   300.000  5000.000 1404.000    21
+1.92317474E+01+1.63154699E-02-5.53448904E-06+8.55059974E-10-4.94583790E-14    2
-1.01971012E+04-7.61674471E+01-4.03105975E+00+7.96101888E-02-7.21655013E-05    3
+3.27610696E-08-5.85584239E-12-3.10973017E+03+4.54324978E+01+0.00000000E+00    4
C6H5OH            L 4/84C   6H   6O   1    0G   300.000  5000.000 1000.        1
+1.49120730E+01+1.83781350E-02-6.19831280E-06+9.19832210E-10-4.92095650E-14    2
-1.83751990E+04-5.59241030E+01-1.69565390E+00+5.22712990E-02-7.20240500E-06    3
-3.58596030E-08+2.04490730E-11-1.32841210E+04+3.25421600E+01-1.15942070E+04    4
C6H5O             T05/02C   6H   5O   1    0G   200.000  6000.000 1000.        1
+1.37221720E+01+1.74688771E-02-6.35504520E-06+1.03492308E-09-6.23410504E-14    2
+2.87274751E+02-4.88181680E+01-4.66204455E-01+4.13443975E-02+1.32412991E-05    3
-5.72872769E-08+2.89763707E-11+4.77858391E+03+2.76990274E+01+6.49467016E+03    4
C6H4OH     4/ 9/ 9 THERMC   6H   5O   1    0G   300.000  5000.000 1402.000    11
+1.73187560E+01+1.36366984E-02-4.68316332E-06+7.29071204E-10-4.23805358E-14    2
+1.14990276E+04-6.89986593E+01-5.99875435E+00+8.59063379E-02-9.12525636E-05    3
+4.72275890E-08-9.35576749E-12+1.78621926E+04+4.99931427E+01+0.00000000E+00    4
OC6H4OH    4/ 9/ 9 THERMC   6H   5O   2    0G   300.000  5000.000 1403.000    11
+2.22718210E+01+1.21038561E-02-4.18429526E-06+6.54475399E-10-3.81746504E-14    2
-2.34827539E+04-9.61035467E+01-8.02205657E+00+1.09403210E-01-1.23489276E-04    3
+6.56286805E-08-1.31527870E-11-1.55949156E+04+5.72175202E+01+0.00000000E+00    4
O-C6H4O2          AK0405C   6H   4O   2    0G   270.000  3000.000 1370.00      1
+1.23614349E+01+2.40491397E-02-1.16529057E-05+2.71332785E-09-2.47593219E-13    2
-1.67079717E+04-4.00310857E+01-2.36179712E+00+6.86058343E-02-6.39129516E-05    3
+3.06903009E-08-5.97357785E-12-1.26704431E+04+3.53724482E+01+0.00000000E+00    4
P-C6H4O2          AK0405C   6H   4O   2    0G   270.000  3000.000 1370.00      1
+1.23423732E+01+2.40612690E-02-1.16565184E-05+2.71393504E-09-2.47643065E-13    2
-2.06185312E+04-4.08244024E+01-2.43170113E+00+6.87937608E-02-6.41382837E-05    3
+3.08126855E-08-5.99832072E-12-1.65696994E+04+3.48309430E+01+0.00000000E+00    4
O-OC6H5OJ  WKM          C   6O   2H   5    0G   300.000  5000.000 1400.000    01
+1.84625733E+01+1.57607263E-02-5.44671499E-06+8.51765760E-10-4.96759541E-14    2
-1.72770226E+02-7.28742484E+01-2.65459198E+00+7.17179095E-02-6.31552372E-05    3
+2.81132946E-08-4.97463333E-12+6.45283150E+03+3.81123139E+01+0.00000000E+00    4
P-OC6H5OJ  WKM          C   6O   2H   5    0G   300.000  5000.000 1400.000    01
+1.82799770E+01+1.59280974E-02-5.50765220E-06+8.61649836E-10-5.02677539E-14    2
-6.25907994E+01-7.25809444E+01-3.29683290E+00+7.27365977E-02-6.36158220E-05    3
+2.80683553E-08-4.92279426E-12+6.73402222E+03+4.09349895E+01+0.00000000E+00    4
P-C6H3O2          AK0505C   6H   3O   2    0G   270.000  3000.000 1290.00      1
+1.22963699E+01+2.15055142E-02-1.07516136E-05+2.57528163E-09-2.41023652E-13    2
+1.15428998E+04-3.72584002E+01-1.57852347E+00+6.55376473E-02-6.50308721E-05    3
+3.32026554E-08-6.86665555E-12+1.51750093E+04+3.31518638E+01+0.00000000E+00    4
C5H6              T 1/90C   5H   6    0    0G   200.000  6000.000 1000.        1
+9.97578480E+00+1.89055430E-02-6.84114610E-06+1.10993400E-09-6.66802360E-14    2
+1.10816930E+04-3.22094540E+01+8.61089570E-01+1.48040310E-02+7.21088950E-05    3
-1.13380550E-07+4.86899720E-11+1.48017550E+04+2.13534530E+01+1.61524850E+04    4
C5H5             TAK0505C   5H   5    0    0G   298.150  3500.000  969.35      1
+1.33675715E+00+3.24793912E-02-1.67587774E-05+4.03514137E-09-3.70739036E-13    2
+3.00730524E+04+1.60315806E+01-3.97555452E+00+7.41370991E-02-1.11803345E-04    3
+9.04628776E-08-2.80999747E-11+3.01769405E+04+3.67153636E+01+0.00000000E+00    4
C5H6-L     2/ 5/ 9 THERMC   5H   6    0    0G   300.000  5000.000 1372.000    21
+1.29600892E+01+1.48953758E-02-5.23622902E-06+8.27916389E-10-4.86464523E-14    2
+2.38180800E+04-4.25312093E+01+3.58448213E+00+3.24459626E-02-1.70150991E-05    3
+4.22715914E-09-4.18452556E-13+2.76514681E+04+9.60644208E+00+0.00000000E+00    4
C#CCVCCJ           GLAR C   5H   5    0    0G   300.000  5000.000 1396.000    11
+1.41230912E+01+1.14233190E-02-3.95851276E-06+6.20128961E-10-3.62097887E-14    2
+4.25158384E+04-5.02942871E+01-6.16143558E-01+5.06466579E-02-4.48561743E-05    3
+2.02459419E-08-3.64542145E-12+4.71532377E+04+2.71623299E+01+0.00000000E+00    4
C5H7       1/22/ 9 WKM  C   5H   7    0    0G   300.000  5000.000 1377.000    31
+1.36630213E+01+1.68061358E-02-5.98746539E-06+9.55341072E-10-5.64951981E-14    2
+1.27238941E+04-5.46331286E+01-6.75118368E+00+6.06461693E-02-4.01260152E-05    3
+1.22051562E-08-1.33459844E-12+2.01365277E+04+5.62694938E+01+0.00000000E+00    4
CVCCJCVC   3/1/95  Z&B  C   5H   7    0    0G   300.000  5000.000 1388.000    21
+1.40879309E+01+1.62398907E-02-5.64768950E-06+8.86857524E-10-5.18698993E-14    2
+1.76798698E+04-5.13735038E+01-2.94595603E+00+5.68783623E-02-4.31336497E-05    3
+1.68169537E-08-2.67926433E-12+2.35156925E+04+3.98188778E+01+0.00000000E+00    4
CVCCVCCJ           Z&B  C   5H   7    0    0G   300.000  5000.000 1386.000    21
+1.47302883E+01+1.59030900E-02-5.57729508E-06+8.80604825E-10-5.16963733E-14    2
+1.74050791E+04-5.42670706E+01-1.60087476E+00+5.38764703E-02-3.96302225E-05    3
+1.49599474E-08-2.31995284E-12+2.31199746E+04+3.35492960E+01+0.00000000E+00    4
CVCCJCVCOH 10/6/95 Z&B  C   5H   7O   1    0G   300.000  5000.000 1397.000    31
+1.67465815E+01+1.58357240E-02-5.44954706E-06+8.49881387E-10-4.94743246E-14    2
-4.30972870E+03-6.19378748E+01-2.91175436E+00+6.69362484E-02-5.71603047E-05    3
+2.48753749E-08-4.33243894E-12+1.96441523E+03+4.17454344E+01+0.00000000E+00    4
CVCCVCCOH  1/23/ 9 WKM  C   5H   8O   1    0G   300.000  5000.000 1396.000    31
+1.63079670E+01+1.79957763E-02-6.03115896E-06+9.23992259E-10-5.31254053E-14    2
-1.58204603E+04-5.84137244E+01-5.31488384E-01+6.06983915E-02-4.81499862E-05    3
+2.00308244E-08-3.38987282E-12-1.03301302E+04+3.07961436E+01+0.00000000E+00    4
C5H5OH     5/ 2/91 THE.MC   5H   6O   1    0G   300.000  5000.000 1398.000    11
+1.53433477E+01+1.50754059E-02-5.13553582E-06+7.95807816E-10-4.61311517E-14    2
-1.19645453E+04-5.85204430E+01-4.26822012E+00+6.62446749E-02-5.68494038E-05    3
+2.46858526E-08-4.26820696E-12-5.75581338E+03+4.47962850E+01+0.00000000E+00    4
C5H5O      5/16/90 THERMC   5H   5O   1    0G   300.000  5000.000 1392.000    01
+1.48322894E+01+1.40483376E-02-4.92302051E-06+7.77041219E-10-4.56103939E-14    2
+1.45523665E+04-5.73228191E+01-2.83112840E+00+5.67277287E-02-4.44757303E-05    3
+1.74924447E-08-2.76004847E-12+2.04992154E+04+3.69634411E+01+0.00000000E+00    4
C5H4OH            T 8/99C   5H   5O   1    0G   200.000  6000.000 1000.        1
+1.33741248E+01+1.51996469E-02-5.45685046E-06+8.80944866E-10-5.27493258E-14    2
+2.20358027E+03-4.59569069E+01-1.28398054E+00+4.90298511E-02-1.35844414E-05    3
-2.92983743E-08+1.90820619E-11+6.37364803E+03+3.08073591E+01+8.00114499E+03    4
C5H4O             T 8/99C   5H   4O   1    0G   200.000  6000.000 1000.        1
+1.00806824E+01+1.61143465E-02-5.83314509E-06+9.46759320E-10-5.68972206E-14    2
+1.94364771E+03-2.94521623E+01+2.64576497E-01+3.34873827E-02+1.67738470E-06    3
-2.96207455E-08+1.54431476E-11+5.11159287E+03+2.35409513E+01+6.64245999E+03    4
C5H3O            TAK0905C   5H   3O   1    0G   300.000  3500.000 1500.00      1
+1.19961781E+01+1.34287065E-02-5.90045309E-06+1.22553862E-09-9.86114716E-14    2
+2.89592010E+04-4.07548249E+01-3.03242604E+00+5.43937201E-02-4.95018348E-05    3
+2.25523751E-08-4.10727920E-12+3.35644081E+04+3.78374823E+01+0.00000000E+00    4
CJVCCVCCVO 2/ 5/ 9 THERMC   5H   5O   1    0G   300.000  5000.000 1396.000    21
+1.62360823E+01+1.18297101E-02-4.11454219E-06+6.46026823E-10-3.77767639E-14    2
+1.93499885E+04-5.83498817E+01-5.06628841E-01+6.04671965E-02-5.97396749E-05    3
+2.96804228E-08-5.76240010E-12+2.42765544E+04+2.82994148E+01+0.00000000E+00    4
CVCCVCCJVO 2/ 5/ 9 THERMC   5H   5O   1    0G   300.000  5000.000 1399.000    11
+1.53178248E+01+1.27352911E-02-4.35882964E-06+6.76912763E-10-3.92771371E-14    2
+7.60582726E+03-5.43599625E+01-2.18492198E-01+5.92100223E-02-5.89241174E-05    3
+2.97411920E-08-5.85244770E-12+1.20600764E+04+2.55968530E+01+0.00000000E+00    4
CJVCCVO    4/ 8/94 THERMC   3H   3O   1    0G   300.000  5000.000 1402.000    11
+1.07482537E+01+6.19822688E-03-2.06130981E-06+3.14418872E-10-1.80309517E-14    2
+1.51410162E+04-3.01266033E+01+1.46654466E+00+3.23390476E-02-3.05588208E-05    3
+1.44081861E-08-2.65600505E-12+1.78850058E+04+1.80850321E+01+0.00000000E+00    4
HOCVCCVO   1/26/ 9 WKM  C   3H   4O   2    0G   300.000  5000.000 1413.000    21
+1.66505478E+01+6.11745137E-03-2.09080785E-06+3.24985683E-10-1.88875073E-14    2
-3.82179939E+04-6.36794754E+01-2.01837189E+00+6.26539783E-02-6.73359280E-05    3
+3.39430425E-08-6.48917648E-12-3.31367523E+04+3.18162860E+01+0.00000000E+00    4
HOCVCCJVO  1/26/ 9 WKM  C   3H   3O   2    0G   300.000  5000.000 1414.000    11
+1.52720985E+01+5.02586331E-03-1.68408578E-06+2.58390706E-10-1.48849424E-14    2
-1.98506828E+04-5.54641734E+01+6.07270082E-01+4.96011303E-02-5.32300885E-05    3
+2.68392951E-08-5.13094510E-12-1.58814562E+04+1.94817133E+01+0.00000000E+00    4
OC5H7O     1/22/ 9 WKM  C   5H   7O   2    0G   300.000  5000.000 1375.000    31
+1.65416953E+01+1.86677673E-02-6.44836048E-06+1.00787611E-09-5.87521858E-14    2
-2.82017168E+04-5.47258181E+01+4.88394767E+00+4.03401300E-02-1.97774150E-05    3
+3.68903501E-09-3.40202384E-14-2.35295942E+04+9.97070337E+00+0.00000000E+00    4
OC4H6O     1/23/ 9 WKM  C   4H   6O   2    0G   300.000  5000.000 1382.000    31
+1.41894774E+01+1.53345510E-02-5.24594862E-06+8.14655154E-10-4.72759368E-14    2
-4.10001835E+04-4.43771751E+01+4.21628848E+00+3.57422725E-02-2.04226185E-05    3
+5.63821367E-09-5.88888993E-13-3.72055911E+04+1.02814620E+01+0.00000000E+00    4
OC4H5O     1/23/ 9 WKM  C   4H   5O   2    0G   300.000  5000.000 1388.000    21
+1.32138775E+01+1.37339051E-02-4.62639517E-06+7.10941370E-10-4.09538499E-14    2
-2.16535271E+04-3.64185255E+01+4.60550978E+00+3.30498712E-02-2.13102363E-05    3
+7.37021089E-09-1.08289438E-12-1.85460831E+04+1.01599453E+01+0.00000000E+00    4
O2CCHOOJ           Z&B  C   2H   1O   4    0G   300.000  5000.000 1682.000    01
+1.09910849E+01+7.46985861E-03-2.75568271E-06+4.51353051E-10-2.72108652E-14    2
-3.51335323E+04-2.11652231E+01+8.91497688E+00+8.60571847E-03+5.24416766E-07    3
-2.79301331E-09+7.62963051E-13-3.40867754E+04-8.72978273E+00+0.00000000E+00    4
C6H5CH3           L 6/87C   7H   8    0    0G   200.000  6000.000 1000.        1
+1.29400340E+01+2.66912870E-02-9.68385050E-06+1.57386290E-09-9.46636010E-14    2
-6.97649080E+02-4.67287850E+01+1.61526630E+00+2.10994380E-02+8.53660180E-05    3
-1.32610660E-07+5.59566040E-11+4.07563000E+03+2.02822100E+01+6.01358350E+03    4
C6H5CH2           IU3/03C  7.H  7.   0.   0.G   250.000  6000.000 1000.        1
+1.47230520E+01+2.30342440E-02-8.48473590E-06+1.39169620E-09-8.42479670E-14    2
+1.79901890E+04-5.59509890E+01-1.23038360E+00+4.89863760E-02+1.38155180E-05    3
-6.25872330E-08+3.15957310E-11+2.31928770E+04+3.05554950E+01+2.50166220E+04    4
C6H4CH3                 C   7H   7    0    0G   300.000  5000.000 1393.000    11
+1.50088040E+01+2.08076711E-02-7.18274868E-06+1.12201995E-09-6.53756838E-14    2
+2.89360689E+04-5.63866198E+01-2.51731357E+00+6.18263711E-02-4.43238513E-05    3
+1.66517959E-08-2.59379321E-12+3.50509401E+04+3.77723973E+01+0.00000000E+00    4
C7H6         G3SX B3LYPTC   7H   6    0    0G   300.000  5000.000 1401.00      1
+1.70564548E+01+1.67766601E-02-5.75637904E-06+8.95748927E-10-5.20574674E-14    2
+3.43929834E+04-6.83510071E+01-3.96406850E+00+7.40750426E-02-6.68009279E-05    3
+3.06821623E-08-5.59258820E-12+4.08575050E+04+4.16088550E+01+0.00000000E+00    4
C7H5         G3SX REF819C   7H   5    0    0G   300.000  5000.000 1404.00      1
+1.65644050E+01+1.44569152E-02-4.91369020E-06+7.59739947E-10-4.39556749E-14    2
+4.96364603E+04-6.29487260E+01-2.77567748E+00+6.97210344E-02-6.63891369E-05    3
+3.18329494E-08-5.98040634E-12+5.53261073E+04+3.73111448E+01+0.00000000E+00    4
BZCOOH                  C   7H   8O   2    0G   300.000  5000.000 1388.000    31
+2.32849942E+01+2.11249905E-02-7.42176803E-06+1.17341778E-09-6.89572814E-14    2
-1.39352842E+04-9.56328725E+01-3.90619768E+00+8.82323518E-02-7.17190897E-05    3
+2.95644635E-08-4.91898930E-12-4.87198921E+03+4.90970451E+01+0.00000000E+00    4
O-O2C6H4CH3  9/21/15    C   7H   7O   2    0G   300.000  5000.000 1408.000    21
+2.12862164E+01+1.93020680E-02-6.48485440E-06+9.95146950E-10-5.72828260E-14    2
+3.19865442E+03-8.60791351E+01-5.17635366E+00+9.32722534E-02-8.64517889E-05    3
+4.02042133E-08-7.33445923E-12+1.10698763E+04+5.15568699E+01+0.00000000E+00    4
OC6H4CH2          012508C   7H   6O   1     G   300.000  5000.000 1000.00      1
+1.24204756E+01+2.70171830E-02-1.09476851E-05+2.02705529E-09-1.40757462E-13    2
+4.49159466E+02-4.10236260E+01-6.21979546E-01+5.14918065E-02-6.11682462E-06    3
-2.88887155E-08+1.45119845E-11+4.44241036E+03+2.88224802E+01+0.00000000E+00    4
C6H5CH2OO  4/10/15      C   7H   7O   2    0G   300.000  5000.000 1390.000    21!HINDER ROTOR NOT CONSIDERED
+2.20121613E+01+2.02138197E-02-7.13572689E-06+1.13165222E-09-6.66401341E-14    2
+4.29764154E+03-9.24408014E+01-4.38932246E+00+8.51137624E-02-6.89728872E-05    3
+2.82508845E-08-4.66501606E-12+1.31191261E+04+4.81693011E+01+0.00000000E+00    4
C6H5CHO    5/16/90 THERMC   7H   6O   1    0G   300.000  5000.000 1386.000    11
+1.74024893E+01+1.89508317E-02-6.58694307E-06+1.03413046E-09-6.04793155E-14    2
-1.31418522E+04-6.83371315E+01-2.37082285E+00+6.28843128E-02-4.26460754E-05    3
+1.39416083E-08-1.74474949E-12-6.11656186E+03+3.85478773E+01+0.00000000E+00    4
C6H5CO                  C   7H   5O   1    0G   300.000  5000.000 1396.000    11
+1.79587471E+01+1.58218495E-02-5.48154854E-06+8.58709339E-10-5.01435299E-14    2
+3.78486787E+03-7.06341032E+01-1.71526142E+00+6.53320500E-02-5.36914036E-05    3
+2.23697440E-08-3.73946626E-12+1.02136508E+04+3.36880709E+01+0.00000000E+00    4
HOC6H4CH3               C   7H   8O   1    0G   300.000  5000.000 1399.000    21
+1.90619388E+01+2.18881056E-02-7.52498751E-06+1.17246043E-09-6.81981400E-14    2
-2.45191428E+04-7.76523319E+01-2.95484914E+00+7.59437004E-02-5.88035350E-05    3
+2.34749185E-08-3.80419645E-12-1.71680056E+04+3.96061710E+01+0.00000000E+00    4
HOC6H4CH2               C   7H   7O   1    0G   300.000  5000.000 1395.000    21
+2.02628865E+01+1.87541796E-02-6.54013354E-06+1.02876061E-09-6.02370606E-14    2
-6.10427929E+03-8.47524281E+01-2.40899264E+00+7.70722558E-02-6.52750566E-05    3
+2.83479112E-08-4.95744925E-12+1.23788601E+03+3.51181131E+01+0.00000000E+00    4
OC6H4CH3                C   7H   7O   1    0G   300.000  5000.000 1392.000    11
+1.81647789E+01+2.08508345E-02-7.23911034E-06+1.13534604E-09-6.63414735E-14    2
-6.88625183E+03-7.15250086E+01-1.85717662E+00+6.67155620E-02-4.70372216E-05    3
+1.67196271E-08-2.39444122E-12+1.36146380E+02+3.62916186E+01+0.00000000E+00    4
OCH3C6H4O  8/ 5/13 THERMC   7H   7O   2    0G   300.000  5000.000 1393.000    11
+2.34089224E+01+1.94710682E-02-6.88461038E-06+1.09305933E-09-6.44198189E-14    2
-2.26138847E+04-1.00700116E+02-7.01264913E+00+9.89740849E-02-8.79431488E-05    3
+3.90945887E-08-6.90477641E-12-1.29339297E+04+5.96245751E+01+0.00000000E+00    4
HOC6H4CH2O              C   7H   7O   2    0G   300.000  5000.000 1372.000    21
+2.19433055E+01+2.04594075E-02-7.26309775E-06+1.15607323E-09-6.82487355E-14    2
-1.66912824E+04-8.93308628E+01+1.68544886E+00+6.20400092E-02-3.79399395E-05    3
+1.06169395E-08-1.05016133E-12-9.04996901E+03+2.15617869E+01+0.00000000E+00    4
HOC6H4CHO               C   7H   6O   2    0G   300.000  5000.000 1398.000    21
+2.21273365E+01+1.63766266E-02-5.56012678E-06+8.60342090E-10-4.98422896E-14    2
-3.66254103E+04-9.10377901E+01-2.48411968E+00+8.02130063E-02-6.92291016E-05    3
+2.97269461E-08-5.04176921E-12-2.88470635E+04+3.86687893E+01+0.00000000E+00    4
HOC6H4CO                C   7H   5O   2    0G   300.000  5000.000 1400.000    21
+2.13743437E+01+1.43756070E-02-4.84732009E-06+7.46563667E-10-4.31103974E-14    2
-1.83638369E+04-8.60689676E+01-7.91109936E-01+7.35177342E-02-6.56772806E-05    3
+2.91823964E-08-5.10216711E-12-1.15203588E+04+3.01664142E+01+0.00000000E+00    4
HOC6H4CH2OOH            C   7H   8O   3    0G   300.000  5000.000 1394.000    41
+2.61613318E+01+2.05361063E-02-7.15910554E-06+1.12622132E-09-6.59585290E-14    2
-3.48441566E+04-1.08404737E+02-2.97566660E+00+9.66654029E-02-8.47224577E-05    3
+3.74478922E-08-6.59470729E-12-2.55751355E+04+4.51493805E+01+0.00000000E+00    4
HOC6H4CH2OO             C   7H   7O   3    0G   300.000  5000.000 1390.000    31
+2.56154733E+01+1.85434725E-02-6.40765412E-06+1.00297172E-09-5.85630540E-14    2
-1.77745474E+04-1.04708103E+02-2.26809341E+00+9.08215743E-02-7.91861666E-05    3
+3.46197851E-08-6.01880047E-12-8.87644654E+03+4.23964585E+01+0.00000000E+00    4
C6H5CH2OH               C   7H   8O   1    0G   300.000  5000.000 1374.000    21
+1.88364511E+01+2.31148752E-02-8.18259004E-06+1.29994648E-09-7.66395338E-14    2
-2.14507156E+04-7.55761963E+01-2.31839760E+00+6.66024713E-02-4.07647160E-05    3
+1.18105957E-08-1.29709981E-12-1.34313628E+04+4.02807703E+01+0.00000000E+00    4
C6H5CHOH                C   7H   7O   1    0G   300.000  5000.000 1369.000    21
+1.87010786E+01+2.07188627E-02-7.36493772E-06+1.17329030E-09-6.93057524E-14    2
+5.13384622E+02-7.34484893E+01-7.47649469E-01+5.95671585E-02-3.49424064E-05    3
+9.19194410E-09-8.16237111E-13+7.99712345E+03+3.34640280E+01+0.00000000E+00    4
C6H5CH2O                C   7H   7O   1    0G   300.000  5000.000 1361.000    11
+1.92483236E+01+2.07494501E-02-7.39239154E-06+1.17943671E-09-6.97421310E-14    2
+5.17232623E+03-7.79664929E+01+2.30480198E-01+5.53611203E-02-2.68816781E-05    3
+3.58435843E-09+4.98228846E-13+1.27838737E+04+2.77013803E+01+0.00000000E+00    4
C6H5C2H5   3/19/ 9 THERMC   8H  10    0    0G   300.000  5000.000 1396.000    21
+2.02158866E+01+2.57181400E-02-8.78778587E-06+1.36387819E-09-7.91252430E-14    2
-6.87601990E+03-8.53188987E+01-5.70126210E+00+8.90606644E-02-6.84365242E-05    3
+2.70624855E-08-4.33907755E-12+1.79229957E+03+5.27926555E+01+0.00000000E+00    4
C6H5CHCH3  4/ 3/ 9 THERMC   8H   9    0    0G   300.000  5000.000 1395.000    11
+2.03767475E+01+2.34923061E-02-8.02742753E-06+1.24595589E-09-7.22895395E-14    2
+1.07287463E+04-8.69308644E+01-3.62245458E+00+8.22327387E-02-6.34562719E-05    3
+2.51893798E-08-4.05353192E-12+1.87480811E+04+4.09318172E+01+0.00000000E+00    4
C6H5CH2CH2 4/ 7/ 9      C   8H   9    0    0G   300.000  5000.000 1397.000    11
+1.97367479E+01+2.34359910E-02-7.88460514E-06+1.21151657E-09-6.98141943E-14    2
+1.82775793E+04-7.90373183E+01-5.03883577E+00+8.49439879E-02-6.65114973E-05    3
+2.66531641E-08-4.29645325E-12+2.64218438E+04+5.25744447E+01+0.00000000E+00    4
C6H5CHOOCH3   3/11 THERMC   8H   9O   2    0G   300.000  5000.000 1391.000    31
+2.39389417E+01+2.55802179E-02-8.93645471E-06+1.40728440E-09-8.24626131E-14    2
-2.90483393E+03-9.84083931E+01-4.15080808E+00+9.63086315E-02-7.90361848E-05    3
+3.37293640E-08-5.86581277E-12+6.40361986E+03+5.07485305E+01+0.00000000E+00    4
C6H5CH2CH2OO  3/11 THERMC   8H   9O   2    0G   300.000  5000.000 1392.000    31
+2.32195676E+01+2.60543894E-02-9.06848696E-06+1.42450939E-09-8.33254784E-14    2
-9.30560896E+02-9.41996431E+01-2.97717571E+00+9.09238597E-02-7.22332479E-05    3
+3.00778320E-08-5.14215828E-12+7.87040761E+03+4.53100220E+01+0.00000000E+00    4
C6H5C2H3          HW /94C   8H   8    0    0G   300.000  3000.000              1
+1.13032130E+01+3.37098870E-02-1.32088850E-05+2.11409620E-09-8.73113770E-14    2
+1.17253880E+04-3.47379190E+01-3.86784930E+00+6.79478650E-02-2.52303330E-05    3
-1.80171450E-08+1.29984700E-11+1.62002690E+04+4.52717700E+01+0.00000000E+00    4
C6H5CCH2   4/ 3/ 9 THERMC   8H   7    0    0G   300.000  5000.000 1387.000    11
+1.92154972E+01+2.02185937E-02-7.07970746E-06+1.11666465E-09-6.55073301E-14    2
+2.44567929E+04-8.09621525E+01-1.75677703E+00+6.93776528E-02-5.15140526E-05    3
+1.96075933E-08-3.05640961E-12+3.17432364E+04+3.16482133E+01+0.00000000E+00    4
C6H5CHCH   4/ 3/ 9 THERMC   8H   7    0    0G   300.000  5000.000 1397.000    11
+1.90927875E+01+1.98909822E-02-6.86981799E-06+1.07370754E-09-6.25902921E-14    2
+3.82661147E+04-7.72000251E+01-3.64383962E+00+7.85604460E-02-6.60358335E-05    3
+2.85738243E-08-4.98068485E-12+4.55975302E+04+4.29246209E+01+0.00000000E+00    4
C14H14 BIBENZYL   T 5/04C 14.H 14.   0.   0.G   200.000  6000.000 1000.        1
+2.65979897E+01+4.68689340E-02-1.69056103E-05+2.73737090E-09-1.64235887E-13    2
+3.18810786E+03-1.14827874E+02+1.30521842E+00+5.76220698E-02+1.22418244E-04    3
-2.18120750E-07+9.59096665E-11+1.26627763E+04+2.90742354E+01+1.63088384E+04    4
C14H13     3/19/ 9 THERMC  14H  13    0    0G   300.000  5000.000 1396.000    21
+3.47417341E+01+3.59337719E-02-1.22450631E-05+1.89794621E-09-1.10038037E-13    2
+1.74795959E+04-1.61420726E+02-9.29192717E+00+1.47032767E-01-1.20211860E-04    3
+4.97625178E-08-8.23851673E-12+3.17775915E+04+7.18644702E+01+0.00000000E+00    4
C14H12     3/19/ 9 THERMC  14H  12    0    0G   300.000  5000.000 1397.000    21
+3.32102692E+01+3.56298722E-02-1.23336159E-05+1.93073037E-09-1.12678018E-13    2
+1.27147671E+04-1.53412616E+02-9.31596441E+00+1.44390141E-01-1.20631407E-04    3
+5.15297757E-08-8.85124801E-12+2.64875194E+04+7.15504888E+01+0.00000000E+00    4
C14H11     3/19/ 9 THERMC  14H  11    0    0G   300.000  5000.000 1395.000    11
+3.27609182E+01+3.39480669E-02-1.17667240E-05+1.84362057E-09-1.07661574E-13    2
+2.92915217E+04-1.51883228E+02-6.70772425E+00+1.32788823E-01-1.07842007E-04    3
+4.47787253E-08-7.50278981E-12+4.22802338E+04+5.76442987E+01+0.00000000E+00    4
C14H13OOH  3/19/ 9 THERMC  14H  14O   2    0G   300.000  5000.000 1395.000    51
+4.01427062E+01+3.93395367E-02-1.37664348E-05+2.17056135E-09-1.27304368E-13    2
-1.39277882E+04-1.84904308E+02-1.04261530E+01+1.68709899E-01-1.42892982E-04    3
+6.15601039E-08-1.06485940E-11+2.47291567E+03+8.26365480E+01+0.00000000E+00    4
C14H13OO   3/19/ 9 THERMC  14H  13O   2    0G   300.000  5000.000 1394.000    41
+3.76701265E+01+3.91886728E-02-1.36838688E-05+2.15430957E-09-1.26216113E-13    2
+4.38748283E+03-1.69872607E+02-9.53800906E+00+1.60095043E-01-1.34982895E-04    3
+5.84090458E-08-1.01919995E-11+1.97390228E+04+7.99308597E+01+0.00000000E+00    4
C14H12OOH  3/19/ 9 THERMC  14H  13O   2    0G   300.000  5000.000 1394.000    41
+4.02968908E+01+3.71210431E-02-1.30088643E-05+2.05309245E-09-1.20495552E-13    2
+3.67900543E+03-1.86479334E+02-8.32529422E+00+1.61762848E-01-1.37724101E-04    3
+5.95672829E-08-1.03363053E-11+1.94259748E+04+7.06782085E+01+0.00000000E+00    4
C14H12O2H-1O2 9/ 9 THERMC  14H  13O   4    0G   300.000  5000.000 1391.000    71
+4.48785960E+01+3.75685709E-02-1.32824040E-05+2.10858085E-09-1.24255944E-13    2
-9.97231472E+03-2.04041648E+02-9.40646930E+00+1.77878119E-01-1.55260847E-04    3
+6.84418245E-08-1.20655066E-11+7.52457116E+03+8.27128410E+01+0.00000000E+00    4
C14H11O-1O2H 19/ 9 THERMC  14H  12O   3    0G   300.000  5000.000 1393.000    41
+4.03057402E+01+3.72594407E-02-1.30902950E-05+2.06942373E-09-1.21596482E-13    2
-2.78034193E+04-1.82398868E+02-7.77794671E+00+1.57347464E-01-1.29564931E-04    3
+5.40605490E-08-9.07699935E-12-1.19364337E+04+7.29984559E+01+0.00000000E+00    4
C14H13O    3/19/ 9 THERMC  14H  13O   1    0G   300.000  5000.000 1397.000    31
+3.62205336E+01+3.75634484E-02-1.29678295E-05+2.02688785E-09-1.18180078E-13    2
+5.74597621E+03-1.65590808E+02-1.19190739E+01+1.59861239E-01-1.33105430E-04    3
+5.60228564E-08-9.42896323E-12+2.13328544E+04+8.92151705E+01+0.00000000E+00    4
C14H12O   10/19/15      C  14H  12O   1    0G   300.000  5000.000 1394.000    31 !USING ANALOGY GROUP TO ESTIMATE
+3.48141204E+01+3.67953648E-02-1.28282619E-05+2.01783856E-09-1.18158524E-13    2
-1.68668837E+04-1.61938007E+02-9.56374055E+00+1.44801295E-01-1.13794706E-04    3
+4.50882665E-08-7.17648586E-12-2.00559523E+03+7.46678724E+01+0.00000000E+00    4
IND       12/16/94 THERMC   9H   8    0     G   300.000  5000.000 1398.000    01
+2.05650080E+01+2.40327712E-02-8.27638045E-06+1.29145387E-09-7.52114721E-14    2
+9.12366072E+03-8.95735971E+01-7.28231243E+00+9.11988088E-02-6.98829415E-05    3
+2.68064158E-08-4.09653374E-12+1.84576190E+04+5.90250983E+01+0.00000000E+00    4
C10H9                   C  10H   90   00    G   300.00   5000.00  1000.00      1
+2.42293900E+01+2.37029600E-02-7.09346000E-06+1.03581400E-09-6.01751500E-14    2
+1.95099300E+04-1.18237400E+02-2.42912400E+00+8.79982900E-02-5.68390900E-05    3
+1.22281800E-08+8.47450100E-13+2.76230400E+04+2.25328200E+01+0.00000000E+00    4
C10H10    11/13/18 THERMC  10H  10O   0    0G   300.000  5000.000 1388.000    01 !UB REFIT 13-11-2018
 2.75025493E+01 2.53421454E-02-8.65098936E-06 1.34348818E-09-7.80290785E-14    2
 1.57619442E+03-1.40866512E+02-4.29107640E+00 9.81011130E-02-6.98930874E-05    3
 2.36467851E-08-3.00135378E-12 1.25239974E+04 3.00159463E+01                   4
C5H5CH3   12/15/94 THERMC   6H   8    0     G   300.000  5000.000 1399.000    11
+1.58460057E+01+2.00902785E-02-6.93497016E-06+1.08339840E-09-6.31318908E-14    2
+3.42821098E+03-6.44405101E+01-6.05214392E+00+7.63737263E-02-6.34619690E-05    3
+2.72515023E-08-4.72538827E-12+1.05143031E+04+5.13368383E+01+0.00000000E+00    4
C9H7  INDENYL     G3B3  H   7C   9O   0N   0G   300.000  3000.000  1000.000    1
+3.65597547E+00+5.74808463E-02-3.42870600E-05+9.70278793E-09-1.05386412E-12    2
+3.06843457E+04+2.57680216E+00-8.73685384E+00+1.03421636E-01-9.23423393E-05    3
+3.75622958E-08-4.40605270E-12+3.31641009E+04+6.28218291E+01+1.95331441E+04    4
C9H6O INDENONE    G3B3  H   6C   9O   1N   0G   300.000  3000.000  1000.000    1
+4.65659248E+00+5.70055822E-02-3.43174199E-05+9.76177442E-09-1.06334037E-12    2
+4.57857140E+03-7.03868477E-01-6.53928778E+00+9.69323286E-02-8.17698656E-05    3
+2.96699474E-08-2.24993392E-12+6.88883578E+03+5.40945996E+01+2.15662372E+04    4
NAPH       2/ 7/95 THERMC  10H   8    0     G   300.000  5000.000 1400.000    01
+2.35897511E+01+2.43823788E-02-8.47570474E-06+1.33051182E-09-7.77992813E-14    2
+6.53423379E+03-1.12133982E+02-8.84119851E+00+1.09328196E-01-9.50844165E-05    3
+4.18320252E-08-7.33414017E-12+1.68163789E+04+5.86791942E+01+0.00000000E+00    4
NAPH-             G3B3  H   7C  10O   0N   0G   300.000  3000.000  1000.000    1
+3.22892303E+00+6.31264486E-02-3.80582381E-05+1.08454069E-08-1.18342512E-12    2
+4.78400840E+04+5.82016697E+00-8.02718034E+00+1.02924518E-01-8.34272010E-05    3
+2.72135383E-08-7.24559554E-13+5.01363344E+04+6.08902264E+01+2.10209869E+04    4
NAPHV             G3B3  H   7C  10O   0N   0G   300.000  3000.000  1000.000    1
+3.29950506E+00+6.30133365E-02-3.79760083E-05+1.08180756E-08-1.18007697E-12    2
+4.76658373E+04+5.41215697E+00-8.00768796E+00+1.03041289E-01-8.38190998E-05    3
+2.76491726E-08-8.88842208E-13+4.99740633E+04+6.07298980E+01+2.10265738E+04    4
NAPHO   THTHOXY   T 7/98C  10H   7O   1    0G   200.000  6000.000  1000.000    1
+2.10591364E+01+2.82563070E-02-1.03328686E-05+1.68867034E-09-1.01974767E-13    2
+4.09143507E+03-8.84963398E+01-1.15176448E+00+6.11354512E-02+3.20151083E-05    3
-9.94285290E-08+4.79990043E-11+1.14058756E+04+3.25584836E+01+1.38887800E+04    4
FLUORENE                C  13H  10          G    300.00   5000.00 1000.00      1
+2.31612871E+01+3.92128530E-02-1.25431510E-05+1.33503890E-09+0.00000000E+00    2
+1.23102892E+04-1.03717257E+02-1.12092800E+01+1.29847800E-01-9.07013380E-05    3
+2.32288460E-08+0.00000000E+00+2.19426600E+04+7.48524200E+01+0.00000000E+00    4
C14H10     3/19/ 9 THERMC  14H  10    0    0G   300.000  5000.000 1387.000    21
+3.35905687E+01+3.03999884E-02-1.05869652E-05+1.66527782E-09-9.75498585E-14    2
+3.04676726E+04-1.56193464E+02-8.67061479E+00+1.30751909E-01-1.00532524E-04    3
+3.78085301E-08-5.59154283E-12+4.47563353E+04+6.98275686E+01+0.00000000E+00    4
C16H10                  C  16H  10          G    300.00   5000.00 1000.00      1
+2.90747022E+01+4.12337670E-02-1.26077060E-05+1.27453580E-09+0.00000000E+00    2
+1.41687238E+04-1.36431347E+02-1.06811200E+01+1.46535400E-01-1.03943520E-04    3
+2.70645390E-08+0.00000000E+00+2.52715000E+04+6.99617500E+01+0.00000000E+00    4
END
